#******
# Preview export LEF
#
#        Preview sub-version 4.4.2.100.41
#
# TECH LIB NAME: tsmc13
#
# RC values have been extracted from TSMC's worst case interconnect
# tables included with CL013G FSG spice model version 1.3P1.
# Document No. T-013-LO-SP-004-PR Rev1.3P1 Jan. 15, 2002
# RC values are also compatible with CL013LV FSG version 1.1
# Document No. T-013-LO-SP-009 Rev1.1 Jan. 29, 2002
#
# Resistance and Capacitance Values
# ---------------------------------
# The LEF technology files included in this directory contain resistance and
# capacitance (RC) values for the purpose of timing driven place & route.
# Please note that the RC values contained in this tech file were created using
# the worst case interconnect models from the foundry and assume a full metal
# route at every grid location on every metal layer, so the values are
# intentionally very conservative. It is assumed that this technology file will
# be used only as a starting point for creating initial timing driven place &
# route runs during the development of your own more accurate RC values,
# tailored to your specific place & route environment. AS A RESULT, TIMING
# NUMBERS DERIVED FROM THESE RC VALUES MAY BE SIGNIFICANTLY SLOWER THAN
# REALITY.
# 
# The RC values used in the LEF technology file are to be used only for timing
# driven place & route. Due to accuracy limitations, please do not attempt to
# use this file for chip-level RC extraction in conjunction with your sign-off
# timing simulations. For chip-level extraction, please use a dedicated
# extraction tool such as HyperExtract, starRC or Simplex, etc.
#
# Antenna Effect Properties
# -------------------------
# Antenna effect properties were modeled based on the following design rule
# document:
#
# Document No. T-013-LO-DR-001 (TSMC 0.13um Logic 1P8M Salicide 1.0V/2.5V,
#                            1.2V/2.5V, 1.0V/3.3V, 1.2V/3.3V Design Rule
#                            version 1.5 8/1/02 )
#
# DO NOT USE SILICON ENSEMBLE OR WROUTE AS A SIGN-OFF VALIDATION FLOW FOR
# PROCESS ANTENNA EFFECT VIOLATIONS.  Foundry DRC command files should always be
# used for sign-off validation of process antenna effect in your design.
#
# $Id: tsmc13fsg_8lm_tech.lef,v 1.3 2004-03-05 19:15:54-08 wching Exp $
#
#******

##############################
# Modified by CIC 2005/07/29 #
##############################
VERSION 5.5 ;
##############################
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

UNITS
    DATABASE MICRONS 2000  ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1

LAYER METAL1
    TYPE ROUTING ;
    WIDTH 0.160 ;
    SPACING 0.180 ;
    SPACING 0.18 LENGTHTHRESHOLD  1.0 ;
    SPACING 0.22 RANGE 0.3 10.0 USELENGTHTHRESHOLD ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.122 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.26 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL1 = 0.117 ohm/sq) = 1.1700e-01
    RESISTANCE RPERSQ      1.1700e-01 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M2-M1-PO1(FOX):0.16:0.18: CAP1 = (Cb_a * PO1(FOX) ratio + Ct_a * M2 ratio) / M1 width = 0.0761773073136342
      # M2-M1-PO1(FOX):0.16:0.18: CAP1 = (6.44e-03 * 1 + 1.11e-02 * 0.401752173913043) / 0.14308 = 0.0761773073136342
      # M3-M1-PO1(FOX):0.16:0.18: CAP2 = (Cb_a * PO1(FOX) ratio + Ct_a * M3 ratio) / M1 width = 0.0163485392787252
      # M3-M1-PO1(FOX):0.16:0.18: CAP2 = (6.44e-03 * 0 + 3.91e-03 * 0.598247826086957) / 0.14308 = 0.0163485392787252
      # CAP = (0.0761773073136342 + 0.0163485392787252) * 0.001 pF/fF = 9.2526e-05
    CAPACITANCE CPERSQDIST 9.2526e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M2-M1-PO1(FOX):0.16:0.18: ECAP1 = Cfb * PO1(FOX) ratio + Cft * M2 ratio = 0.019456896
      # M2-M1-PO1(FOX):0.16:0.18: ECAP1 = 1.65e-02 * 1 + 7.36e-03 * 0.401752173913043 = 0.019456896
      # M3-M1-PO1(FOX):0.16:0.18: ECAP2 = Cfb * PO1(FOX) ratio + Cft * M3 ratio = 0.00176483108695652
      # M3-M1-PO1(FOX):0.16:0.18: ECAP2 = 1.71e-02 * 0 + 2.95e-03 * 0.598247826086957 = 0.00176483108695652
      # M3-M1-PO1(FOX):0.16:0.18: Cc = 7.88e-02
      # ECAP = (0.019456896 + 0.00176483108695652 + 7.88e-02) * 0.001 pF/fF = 1.0002e-04
    EDGECAPACITANCE        1.0002e-04 ;
END METAL1

LAYER VIA12
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA12

LAYER METAL2
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL2 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M3-M2-M1:0.2:0.21: CAP1 = (Cb_a * M1 ratio + Ct_a * M3 ratio) / M2 width = 0.073567268827456
      # M3-M2-M1:0.2:0.21: CAP1 = (1.43e-02 * 0.5 + 1.43e-02 * 0.450746341463415) / 0.184806 = 0.073567268827456
      # M4-M2-PO1(FOX):0.2:0.21: CAP2 = (Cb_a * PO1(FOX) ratio + Ct_a * M4 ratio) / M2 width = 0.03232433457577
      # M4-M2-PO1(FOX):0.2:0.21: CAP2 = (6.40e-03 * 0.5 + 5.05e-03 * 0.549253658536585) / 0.184806 = 0.03232433457577
      # CAP = (0.073567268827456 + 0.03232433457577) * 0.001 pF/fF = 1.0589e-04
    CAPACITANCE CPERSQDIST 1.0589e-04 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M3-M2-M1:0.2:0.21: ECAP1 = Cfb * M1 ratio + Cft * M3 ratio = 0.00782774687804878
      # M3-M2-M1:0.2:0.21: ECAP1 = 8.11e-03 * 0.5 + 8.37e-03 * 0.450746341463415 = 0.00782774687804878
      # M4-M2-PO1(FOX):0.2:0.21: ECAP2 = Cfb * PO1(FOX) ratio + Cft * M4 ratio = 0.00411886541463415
      # M4-M2-PO1(FOX):0.2:0.21: ECAP2 = 4.36e-03 * 0.5 + 3.53e-03 * 0.549253658536585 = 0.00411886541463415
      # M4-M2-PO1(FOX):0.2:0.21: Cc = 8.65e-02
      # ECAP = (0.00782774687804878 + 0.00411886541463415 + 8.65e-02) * 0.001 pF/fF = 9.8447e-05
    EDGECAPACITANCE        9.8447e-05 ;
END METAL2

LAYER VIA23
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA23

LAYER METAL3
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL3 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M4-M3-M2:0.2:0.21: CAP1 = (Cb_a * M2 ratio + Ct_a * M4 ratio) / M3 width = 0.0621739130434783
      # M4-M3-M2:0.2:0.21: CAP1 = (1.43e-02 * 0.401752173913043 + 1.43e-02 * 0.401752173913043) / 0.184806 = 0.0621739130434783
      # M5-M3-M1:0.2:0.21: CAP2 = (Cb_a * M1 ratio + Ct_a * M5 ratio) / M3 width = 0.0326953835020414
      # M5-M3-M1:0.2:0.21: CAP2 = (5.05e-03 * 0.598247826086957 + 5.05e-03 * 0.598247826086957) / 0.184806 = 0.0326953835020414
      # CAP = (0.0621739130434783 + 0.0326953835020414) * 0.001 pF/fF = 9.4869e-05
    CAPACITANCE CPERSQDIST 9.4869e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M4-M3-M2:0.2:0.21: ECAP1 = Cfb * M2 ratio + Cft * M4 ratio = 0.00662087582608696
      # M4-M3-M2:0.2:0.21: ECAP1 = 8.11e-03 * 0.401752173913043 + 8.37e-03 * 0.401752173913043 = 0.00662087582608696
      # M5-M3-M1:0.2:0.21: ECAP2 = Cfb * M1 ratio + Cft * M5 ratio = 0.00433729673913043
      # M5-M3-M1:0.2:0.21: ECAP2 = 3.63e-03 * 0.598247826086957 + 3.62e-03 * 0.598247826086957 = 0.00433729673913043
      # M5-M3-M1:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00662087582608696 + 0.00433729673913043 + 8.70e-02) * 0.001 pF/fF = 9.7958e-05
    EDGECAPACITANCE        9.7958e-05 ;
END METAL3

LAYER VIA34
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA34

LAYER METAL4
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL4 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M5-M4-M3:0.2:0.21: CAP1 = (Cb_a * M3 ratio + Ct_a * M5 ratio) / M4 width = 0.0697560975609756
      # M5-M4-M3:0.2:0.21: CAP1 = (1.43e-02 * 0.450746341463415 + 1.43e-02 * 0.450746341463415) / 0.184806 = 0.0697560975609756
      # M6-M4-M2:0.2:0.21: CAP2 = (Cb_a * M2 ratio + Ct_a * M6 ratio) / M4 width = 0.0300177588997084
      # M6-M4-M2:0.2:0.21: CAP2 = (5.05e-03 * 0.549253658536585 + 5.05e-03 * 0.549253658536585) / 0.184806 = 0.0300177588997084
      # CAP = (0.0697560975609756 + 0.0300177588997084) * 0.001 pF/fF = 9.9774e-05
    CAPACITANCE CPERSQDIST 9.9774e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M5-M4-M3:0.2:0.21: ECAP1 = Cfb * M3 ratio + Cft * M5 ratio = 0.00742829970731707
      # M5-M4-M3:0.2:0.21: ECAP1 = 8.11e-03 * 0.450746341463415 + 8.37e-03 * 0.450746341463415 = 0.00742829970731707
      # M6-M4-M2:0.2:0.21: ECAP2 = Cfb * M2 ratio + Cft * M6 ratio = 0.00398208902439024
      # M6-M4-M2:0.2:0.21: ECAP2 = 3.63e-03 * 0.549253658536585 + 3.62e-03 * 0.549253658536585 = 0.00398208902439024
      # M6-M4-M2:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00742829970731707 + 0.00398208902439024 + 8.70e-02) * 0.001 pF/fF = 9.8410e-05
    EDGECAPACITANCE        9.8410e-05 ;
END METAL4

LAYER VIA45
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA45

LAYER METAL5
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.410 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL5 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M6-M5-M4:0.2:0.21: CAP1 = (Cb_a * M4 ratio + Ct_a * M6 ratio) / M5 width = 0.0621739130434783
      # M6-M5-M4:0.2:0.21: CAP1 = (1.43e-02 * 0.401752173913043 + 1.43e-02 * 0.401752173913043) / 0.184806 = 0.0621739130434783
      # M7-M5-M3:0.2:0.21: CAP2 = (Cb_a * M3 ratio + Ct_a * M7 ratio) / M5 width = 0.0326953835020414
      # M7-M5-M3:0.2:0.21: CAP2 = (5.05e-03 * 0.598247826086957 + 5.05e-03 * 0.598247826086957) / 0.184806 = 0.0326953835020414
      # CAP = (0.0621739130434783 + 0.0326953835020414) * 0.001 pF/fF = 9.4869e-05
    CAPACITANCE CPERSQDIST 9.4869e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M6-M5-M4:0.2:0.21: ECAP1 = Cfb * M4 ratio + Cft * M6 ratio = 0.00662087582608696
      # M6-M5-M4:0.2:0.21: ECAP1 = 8.11e-03 * 0.401752173913043 + 8.37e-03 * 0.401752173913043 = 0.00662087582608696
      # M7-M5-M3:0.2:0.21: ECAP2 = Cfb * M3 ratio + Cft * M7 ratio = 0.00433729673913043
      # M7-M5-M3:0.2:0.21: ECAP2 = 3.63e-03 * 0.598247826086957 + 3.62e-03 * 0.598247826086957 = 0.00433729673913043
      # M7-M5-M3:0.2:0.21: Cc = 8.70e-02
      # ECAP = (0.00662087582608696 + 0.00433729673913043 + 8.70e-02) * 0.001 pF/fF = 9.7958e-05
    EDGECAPACITANCE        9.7958e-05 ;
END METAL5

LAYER VIA56
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA56

LAYER METAL6
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.460 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL6 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M7-M6-M5:0.2:0.21: CAP1 = (Cb_a * M5 ratio + Ct_a * M7 ratio) / M6 width = 0.058130081300813
      # M7-M6-M5:0.2:0.21: CAP1 = (1.43e-02 * 0.450746341463415 + 1.43e-02 * 0.30049756097561) / 0.184806 = 0.058130081300813
      # M8-M6-M4:0.2:0.21: CAP2 = (Cb_a * M4 ratio + Ct_a * M8 ratio) / M6 width = 0.0322687688579428
      # M8-M6-M4:0.2:0.21: CAP2 = (5.05e-03 * 0.549253658536585 + 4.56e-03 * 0.69950243902439) / 0.184806 = 0.0322687688579428
      # CAP = (0.058130081300813 + 0.0322687688579428) * 0.001 pF/fF = 9.0399e-05
    CAPACITANCE CPERSQDIST 9.0399e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M7-M6-M5:0.2:0.21: ECAP1 = Cfb * M5 ratio + Cft * M7 ratio = 0.00617071741463415
      # M7-M6-M5:0.2:0.21: ECAP1 = 8.11e-03 * 0.450746341463415 + 8.37e-03 * 0.30049756097561 = 0.00617071741463415
      # M8-M6-M4:0.2:0.21: ECAP2 = Cfb * M4 ratio + Cft * M8 ratio = 0.00442002941463415
      # M8-M6-M4:0.2:0.21: ECAP2 = 3.73e-03 * 0.549253658536585 + 3.39e-03 * 0.69950243902439 = 0.00442002941463415
      # M8-M6-M4:0.2:0.21: Cc = 8.73e-02
      # ECAP = (0.00617071741463415 + 0.00442002941463415 + 8.73e-02) * 0.001 pF/fF = 9.7891e-05
    EDGECAPACITANCE        9.7891e-05 ;
END METAL6

LAYER VIA67
    TYPE CUT ;
    SPACING 0.220 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA67

LAYER METAL7
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.210 ;
    SPACING 0.24 RANGE 0.39 10.0 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 0.615 ;
    OFFSET 0.205 ;
    DIRECTION HORIZONTAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.144 ;
    MINIMUMCUT 2 WIDTH 1.40 ;
    THICKNESS 0.35 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 43062 ) ( 1 43436 ) ) ;
      # (Worst case resistance model for METAL7 = 0.077 ohm/sq) = 7.7000e-02
    RESISTANCE RPERSQ      7.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M8-M7-M6:0.2:0.41: CAP1 = (Cb_a * M6 ratio + Ct_a * M8 ratio) / M7 width = 0.0521304244309779
      # M8-M7-M6:0.2:0.41: CAP1 = (1.43e-02 * 0.401752173913043 + 1.10e-02 * 0.353541739130435) / 0.184806 = 0.0521304244309779
      # M7-M5:0.2:0.41: CAP2 = Ca * M5 ratio / M7 width = 0.0163476917510207
      # M7-M5:0.2:0.41: CAP2 = 5.05e-03 * 0.598247826086957 / 0.184806 = 0.0163476917510207
      # CAP = (0.0521304244309779 + 0.0163476917510207) * 0.001 pF/fF = 6.8478e-05
    CAPACITANCE CPERSQDIST 6.8478e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M8-M7-M6:0.2:0.41: ECAP1 = Cfb * M6 ratio + Cft * M8 ratio = 0.00965490626086957
      # M8-M7-M6:0.2:0.41: ECAP1 = 1.40e-02 * 0.401752173913043 + 1.14e-02 * 0.353541739130435 = 0.00965490626086957
      # M7-M5:0.2:0.41: ECAP2 = Cf * M5 ratio = 0.00506715908695652
      # M7-M5:0.2:0.41: ECAP2 = 8.47e-03 * 0.598247826086957 = 0.00506715908695652
      # M7-M5:0.2:0.41: Cc = 5.33e-02
      # ECAP = (0.00965490626086957 + 0.00506715908695652 + 5.33e-02) * 0.001 pF/fF = 6.8022e-05
    EDGECAPACITANCE        6.8022e-05 ;
END METAL7

LAYER VIA78
    TYPE CUT ;
    SPACING 0.350 ;
    ANTENNAAREARATIO 50 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 50 ) ( 0.159 50 ) ( 0.16 933 ) ( 1 1110 ) ) ;
END VIA78

LAYER METAL8
    TYPE ROUTING ;
    WIDTH 0.440 ;
    SPACING 0.460 ;
    SPACING 0.60 RANGE 10.05 100000.0 ;
    PITCH 1.150 ;
    OFFSET 0.230 ;
    DIRECTION VERTICAL ;
##############################
# Modified by CIC 2005/07/29 #
##############################
    MAXWIDTH 11.0 ;
##############################
    AREA 0.562 ;
    MINIMUMCUT 2 WIDTH 1.80 ;
    THICKNESS 0.90 ;
    ANTENNACUMAREARATIO 5496 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5496 ) ( 0.159 5496 ) ( 0.16 51270 ) ( 1 57980 ) ) ;
      # (Worst case resistance model for METAL8 = 0.027 ohm/sq) = 2.7000e-02
    RESISTANCE RPERSQ      2.7000e-02 ;
      # CAP = (CAP1 + CAP2) * 0.001 pF/fF
      # M8-M7:0.44:0.66: CAP1 = Ca * M7 ratio / M8 width = 0.0178861876602966
      # M8-M7:0.44:0.66: CAP1 = 2.42e-02 * 0.30049756097561 / 0.406573 = 0.0178861876602966
      # M8-M6:0.44:0.66: CAP2 = Ca * M6 ratio / M8 width = 0.0172048424028253
      # M8-M6:0.44:0.66: CAP2 = 1.00e-02 * 0.69950243902439 / 0.406573 = 0.0172048424028253
      # CAP = (0.0178861876602966 + 0.0172048424028253) * 0.001 pF/fF = 3.5091e-05
    CAPACITANCE CPERSQDIST 3.5091e-05 ;
      # ECAP = (ECAP1 + ECAP2 + Cc) * 0.001 pF/fF
      # M8-M7:0.44:0.66: ECAP1 = Cf * M7 ratio = 0.00558925463414634
      # M8-M7:0.44:0.66: ECAP1 = 1.86e-02 * 0.30049756097561 = 0.00558925463414634
      # M8-M6:0.44:0.66: ECAP2 = Cf * M6 ratio = 0.00647739258536585
      # M8-M6:0.44:0.66: ECAP2 = 9.26e-03 * 0.69950243902439 = 0.00647739258536585
      # M8-M6:0.44:0.66: Cc = 7.25e-02
      # ECAP = (0.00558925463414634 + 0.00647739258536585 + 7.25e-02) * 0.001 pF/fF = 8.4567e-05
    EDGECAPACITANCE        8.4567e-05 ;
END METAL8

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIARULE VIA1ARRAY GENERATE
    LAYER METAL1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA1ARRAY

VIARULE VIA2ARRAY GENERATE
    LAYER METAL2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA2ARRAY

VIARULE VIA3ARRAY GENERATE
    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA3ARRAY

VIARULE VIA4ARRAY GENERATE
    LAYER METAL4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA4ARRAY

VIARULE VIA5ARRAY GENERATE
    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA5ARRAY

VIARULE VIA6ARRAY GENERATE
    LAYER METAL6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        SPACING 0.480 BY 0.480 ;
END VIA6ARRAY

VIARULE VIA7ARRAY GENERATE
    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.050 ;
        METALOVERHANG 0.000 ;

    LAYER METAL8 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER VIA78 ;
        RECT -0.180 -0.180 0.180 0.180 ;
        SPACING 0.900 BY 0.900 ;
END VIA7ARRAY

VIARULE TURNM1 GENERATE
    LAYER METAL1 ;
        DIRECTION VERTICAL ;

    LAYER METAL1 ;
        DIRECTION HORIZONTAL ;
END TURNM1

VIARULE TURNM2 GENERATE
    LAYER METAL2 ;
        DIRECTION VERTICAL ;

    LAYER METAL2 ;
        DIRECTION HORIZONTAL ;
END TURNM2

VIARULE TURNM3 GENERATE
    LAYER METAL3 ;
        DIRECTION VERTICAL ;

    LAYER METAL3 ;
        DIRECTION HORIZONTAL ;
END TURNM3

VIARULE TURNM4 GENERATE
    LAYER METAL4 ;
        DIRECTION VERTICAL ;

    LAYER METAL4 ;
        DIRECTION HORIZONTAL ;
END TURNM4

VIARULE TURNM5 GENERATE
    LAYER METAL5 ;
        DIRECTION VERTICAL ;

    LAYER METAL5 ;
        DIRECTION HORIZONTAL ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER METAL6 ;
        DIRECTION VERTICAL ;

    LAYER METAL6 ;
        DIRECTION HORIZONTAL ;
END TURNM6

VIARULE TURNM7 GENERATE
    LAYER METAL7 ;
        DIRECTION VERTICAL ;

    LAYER METAL7 ;
        DIRECTION HORIZONTAL ;
END TURNM7

VIARULE TURNM8 GENERATE
    LAYER METAL8 ;
        DIRECTION VERTICAL ;

    LAYER METAL8 ;
        DIRECTION HORIZONTAL ;
END TURNM8

SPACING
    SAMENET METAL1 METAL1 0.180  ;
    SAMENET METAL2 METAL2 0.210  STACK ;
    SAMENET METAL3 METAL3 0.210  STACK ;
    SAMENET METAL4 METAL4 0.210  STACK ;
    SAMENET METAL5 METAL5 0.210  STACK ;
    SAMENET METAL6 METAL6 0.210  STACK ;
    SAMENET METAL7 METAL7 0.210  STACK ;
    SAMENET METAL8 METAL8 0.460  ;
    SAMENET VIA12 VIA12 0.220  ;
    SAMENET VIA23 VIA23 0.220  ;
    SAMENET VIA34 VIA34 0.220  ;
    SAMENET VIA45 VIA45 0.220  ;
    SAMENET VIA56 VIA56 0.220  ;
    SAMENET VIA67 VIA67 0.220  ;
    SAMENET VIA78 VIA78 0.350  ;
    SAMENET VIA12 VIA23 0.0 STACK ;
    SAMENET VIA23 VIA34 0.0 STACK ;
    SAMENET VIA34 VIA45 0.0 STACK ;
    SAMENET VIA45 VIA56 0.0 STACK ;
    SAMENET VIA56 VIA67 0.0 STACK ;
    SAMENET VIA67 VIA78 0.0 STACK ;
END SPACING

VIA VIA12_H DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA12_H

VIA VIA12_V DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA12_V

VIA VIA12_X DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA12_X

VIA VIA12_XR DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA12_XR

VIA VIA23_H DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA23_H

VIA VIA23_V DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_V

VIA VIA23_X DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_X

VIA VIA23_XR DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA23_XR

VIA VIA34_H DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA34_H

VIA VIA34_V DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_V

VIA VIA34_X DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_X

VIA VIA34_XR DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA34_XR

VIA VIA45_H DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA45_H

VIA VIA45_V DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_V

VIA VIA45_X DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_X

VIA VIA45_XR DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA45_XR

VIA VIA56_H DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA56_H

VIA VIA56_V DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_V

VIA VIA56_X DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_X

VIA VIA56_XR DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA56_XR

VIA VIA67_H DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA67_H

VIA VIA67_V DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_V

VIA VIA67_X DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_X

VIA VIA67_XR DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA67_XR

VIA VIA78_H DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.23 -0.19 0.23 0.19 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_H

VIA VIA78_V DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_V

VIA VIA78_XR DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 6.3000e-01
    RESISTANCE 6.3000e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 0.27 ;
END VIA78_XR

VIA VIA23_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL2 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA23_TOS

VIA VIA34_TOS_E DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.580 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_TOS_E

VIA VIA34_TOS_W DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL3 ;
        RECT -0.580 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA34_TOS_W

VIA VIA45_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL4 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA45_TOS

VIA VIA56_TOS_E DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.580 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_TOS_E

VIA VIA56_TOS_W DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL5 ;
        RECT -0.580 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.145 ;
END VIA56_TOS_W

VIA VIA67_TOS DEFAULT TOPOFSTACKONLY
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 1.0200e+00
    RESISTANCE 1.0200e+00 ;
    LAYER METAL6 ;
        RECT -0.1 -0.370 0.1 0.370 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.145 0.1 ;
END VIA67_TOS

VIA VIA12_2CUT_E DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.145 -0.105 0.625 0.105 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA12_2CUT_E

VIA VIA12_2CUT_W DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.625 -0.105 0.145 0.105 ;
    LAYER VIA12 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA12_2CUT_W

VIA VIA12_2CUT_N DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.105 -0.145 0.105 0.625 ;
    LAYER VIA12 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA12_2CUT_N

VIA VIA12_2CUT_S DEFAULT
      # (Worst case resistance model for VIA12 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL1 ;
        RECT -0.105 -0.625 0.105 0.145 ;
    LAYER VIA12 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL2 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA12_2CUT_S

VIA VIA23_2CUT_E DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA23_2CUT_E

VIA VIA23_2CUT_W DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA23 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA23_2CUT_W

VIA VIA23_2CUT_N DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA23 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA23_2CUT_N

VIA VIA23_2CUT_S DEFAULT
      # (Worst case resistance model for VIA23 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL2 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA23 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL3 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA23_2CUT_S

VIA VIA34_2CUT_E DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA34_2CUT_E

VIA VIA34_2CUT_W DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA34 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA34_2CUT_W

VIA VIA34_2CUT_N DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA34 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA34_2CUT_N

VIA VIA34_2CUT_S DEFAULT
      # (Worst case resistance model for VIA34 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL3 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA34 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL4 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA34_2CUT_S

VIA VIA45_2CUT_E DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA45_2CUT_E

VIA VIA45_2CUT_W DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA45 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA45_2CUT_W

VIA VIA45_2CUT_N DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA45 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA45_2CUT_N

VIA VIA45_2CUT_S DEFAULT
      # (Worst case resistance model for VIA45 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL4 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA45 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL5 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA45_2CUT_S

VIA VIA56_2CUT_E DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA56_2CUT_E

VIA VIA56_2CUT_W DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA56 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA56_2CUT_W

VIA VIA56_2CUT_N DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA56 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA56_2CUT_N

VIA VIA56_2CUT_S DEFAULT
      # (Worst case resistance model for VIA56 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL5 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA56 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL6 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA56_2CUT_S

VIA VIA67_2CUT_E DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.145 -0.1 0.625 0.1 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT 0.385 -0.095 0.575 0.095 ;
    LAYER METAL7 ;
        RECT -0.145 -0.1 0.625 0.1 ;
END VIA67_2CUT_E

VIA VIA67_2CUT_W DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.625 -0.1 0.145 0.1 ;
    LAYER VIA67 ;
        RECT -0.575 -0.095 -0.385 0.095 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.625 -0.1 0.145 0.1 ;
END VIA67_2CUT_W

VIA VIA67_2CUT_N DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.1 -0.145 0.1 0.625 ;
    LAYER VIA67 ;
        RECT -0.095 -0.095 0.095 0.095 ;
        RECT -0.095 0.385 0.095 0.575 ;
    LAYER METAL7 ;
        RECT -0.1 -0.145 0.1 0.625 ;
END VIA67_2CUT_N

VIA VIA67_2CUT_S DEFAULT
      # (Worst case resistance model for VIA67 = 1.02 ohm/ct) = 5.1000e-01
    RESISTANCE 5.1000e-01 ;
    LAYER METAL6 ;
        RECT -0.1 -0.625 0.1 0.145 ;
    LAYER VIA67 ;
        RECT -0.095 -0.575 0.095 -0.385 ;
        RECT -0.095 -0.095 0.095 0.095 ;
    LAYER METAL7 ;
        RECT -0.1 -0.625 0.1 0.145 ;
END VIA67_2CUT_S

VIA VIA78_2CUT_E DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.23 -0.19 1.13 0.19 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT 0.72 -0.18 1.08 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 1.17 0.27 ;
END VIA78_2CUT_E

VIA VIA78_2CUT_W DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -1.13 -0.19 0.23 0.19 ;
    LAYER VIA78 ;
        RECT -1.08 -0.18 -0.72 0.18 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -1.17 -0.27 0.27 0.27 ;
END VIA78_2CUT_W

VIA VIA78_2CUT_N DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -0.23 0.19 1.13 ;
    LAYER VIA78 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        RECT -0.18 0.72 0.18 1.08 ;
    LAYER METAL8 ;
        RECT -0.27 -0.27 0.27 1.17 ;
END VIA78_2CUT_N

VIA VIA78_2CUT_S DEFAULT
      # (Worst case resistance model for VIA78 = 0.63 ohm/ct) = 3.1500e-01
    RESISTANCE 3.1500e-01 ;
    LAYER METAL7 ;
        RECT -0.19 -1.13 0.19 0.23 ;
    LAYER VIA78 ;
        RECT -0.18 -1.08 0.18 -0.72 ;
        RECT -0.18 -0.18 0.18 0.18 ;
    LAYER METAL8 ;
        RECT -0.27 -1.17 0.27 0.27 ;
END VIA78_2CUT_S

SITE TSM13SITE
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.460 BY 3.690 ;
END TSM13SITE

MACRO FILL64
    CLASS CORE SPACER ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 29.440 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 29.440 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 29.440 3.940 ;
        END
    END VDD
END FILL64

MACRO FILL32
    CLASS CORE SPACER ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 14.720 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 14.720 3.940 ;
        END
    END VDD
END FILL32

MACRO FILL16
    CLASS CORE SPACER ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 7.360 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 7.360 3.940 ;
        END
    END VDD
END FILL16

MACRO FILL8
    CLASS CORE SPACER ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 3.680 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 3.680 3.940 ;
        END
    END VDD
END FILL8

MACRO FILL4
    CLASS CORE SPACER ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.840 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 1.840 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 1.840 3.940 ;
        END
    END VDD
END FILL4

MACRO FILL2
    CLASS CORE SPACER ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.920 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.920 3.940 ;
        END
    END VDD
END FILL2

MACRO FILL1
    CLASS CORE SPACER ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.460 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.460 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.460 3.940 ;
        END
    END VDD
END FILL1

MACRO ANTENNA
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 0.875 0.590 2.385 ;
        RECT  0.125 0.875 0.330 1.185 ;
        END
        ANTENNADIFFAREA     1.4270 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.250 0.920 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.440 0.920 3.940 ;
        END
    END VDD
END ANTENNA

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.105 0.795 1.580 ;
        RECT  0.585 1.035 0.785 1.580 ;
        RECT  0.525 1.035 0.585 1.355 ;
        END
        ANTENNADIFFAREA     0.1428 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 -0.250 0.920 0.250 ;
        RECT  0.125 -0.250 0.725 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 3.440 0.920 3.940 ;
        RECT  0.315 2.700 0.575 3.940 ;
        RECT  0.000 3.440 0.315 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.315 1.760 0.575 2.390 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.920 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 2.110 0.795 2.400 ;
        RECT  0.525 1.955 0.785 2.555 ;
        END
        ANTENNADIFFAREA     0.2176 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 -0.250 0.920 0.250 ;
        RECT  0.385 -0.250 0.645 0.405 ;
        RECT  0.000 -0.250 0.385 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 3.440 0.920 3.940 ;
        RECT  0.125 2.875 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.545 1.035 0.645 1.295 ;
        RECT  0.385 1.035 0.545 1.675 ;
        RECT  0.125 1.515 0.385 1.775 ;
    END
END TIEHI

MACRO DLY4X4
    CLASS CORE ;
    FOREIGN DLY4X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY4X4

MACRO DLY3X4
    CLASS CORE ;
    FOREIGN DLY3X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY3X4

MACRO DLY2X4
    CLASS CORE ;
    FOREIGN DLY2X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY2X4

MACRO DLY1X4
    CLASS CORE ;
    FOREIGN DLY1X4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.140 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.105 4.015 1.990 ;
        RECT  3.830 1.005 4.005 1.990 ;
        RECT  3.805 0.880 3.830 1.990 ;
        RECT  3.745 0.880 3.805 1.205 ;
        RECT  3.575 1.790 3.805 1.990 ;
        RECT  3.485 0.605 3.745 1.205 ;
        RECT  3.505 1.790 3.575 2.605 ;
        RECT  3.375 1.790 3.505 3.005 ;
        RECT  3.345 2.335 3.375 3.005 ;
        RECT  3.245 2.405 3.345 3.005 ;
        END
        ANTENNADIFFAREA     0.7788 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.295 1.590 0.795 1.990 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 -0.250 4.140 0.250 ;
        RECT  2.975 -0.250 3.235 1.075 ;
        RECT  0.785 -0.250 2.975 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 3.440 4.140 3.940 ;
        RECT  3.755 2.255 4.015 3.940 ;
        RECT  2.955 3.440 3.755 3.940 ;
        RECT  2.695 3.285 2.955 3.940 ;
        RECT  0.785 3.440 2.695 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.585 3.195 1.845 ;
        RECT  2.935 1.255 3.095 2.220 ;
        RECT  2.155 1.255 2.935 1.415 ;
        RECT  2.155 2.060 2.935 2.220 ;
        RECT  2.275 1.595 2.535 1.855 ;
        RECT  1.725 1.645 2.275 1.805 ;
        RECT  1.995 1.035 2.155 1.415 ;
        RECT  1.995 2.060 2.155 2.770 ;
        RECT  1.895 1.035 1.995 1.295 ;
        RECT  1.895 2.510 1.995 2.770 ;
        RECT  1.715 0.525 1.755 0.785 ;
        RECT  1.715 1.645 1.725 2.260 ;
        RECT  1.555 0.525 1.715 2.260 ;
        RECT  1.495 0.525 1.555 0.785 ;
        RECT  1.465 2.000 1.555 2.260 ;
        RECT  1.135 1.495 1.235 1.755 ;
        RECT  0.975 1.245 1.135 2.330 ;
        RECT  0.385 1.245 0.975 1.405 ;
        RECT  0.385 2.170 0.975 2.330 ;
        RECT  0.125 1.035 0.385 1.405 ;
        RECT  0.125 2.170 0.385 2.770 ;
    END
END DLY1X4

MACRO DLY4X1
    CLASS CORE ;
    FOREIGN DLY4X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY4X1

MACRO DLY3X1
    CLASS CORE ;
    FOREIGN DLY3X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY3X1

MACRO DLY2X1
    CLASS CORE ;
    FOREIGN DLY2X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY2X1

MACRO DLY1X1
    CLASS CORE ;
    FOREIGN DLY1X1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 1.035 3.555 2.555 ;
        RECT  3.370 1.035 3.395 1.355 ;
        RECT  3.370 1.925 3.395 2.555 ;
        RECT  3.295 1.035 3.370 1.295 ;
        RECT  3.295 1.955 3.370 2.555 ;
        END
        ANTENNADIFFAREA     0.3306 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.245 0.795 1.665 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 -0.250 3.680 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  0.785 -0.250 2.835 0.250 ;
        RECT  0.525 -0.250 0.785 0.405 ;
        RECT  0.000 -0.250 0.525 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 3.440 3.680 3.940 ;
        RECT  2.835 3.285 3.095 3.940 ;
        RECT  0.785 3.440 2.835 3.940 ;
        RECT  0.525 3.285 0.785 3.940 ;
        RECT  0.000 3.440 0.525 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 1.515 3.195 1.775 ;
        RECT  2.935 1.020 3.095 2.115 ;
        RECT  2.125 1.020 2.935 1.180 ;
        RECT  2.155 1.955 2.935 2.115 ;
        RECT  2.345 1.470 2.605 1.730 ;
        RECT  1.725 1.520 2.345 1.680 ;
        RECT  1.995 1.955 2.155 2.785 ;
        RECT  1.965 0.525 2.125 1.180 ;
        RECT  1.895 2.525 1.995 2.785 ;
        RECT  1.865 0.525 1.965 0.785 ;
        RECT  1.565 1.035 1.725 2.275 ;
        RECT  1.465 1.035 1.565 1.295 ;
        RECT  1.465 2.015 1.565 2.275 ;
        RECT  1.015 1.595 1.265 2.005 ;
        RECT  0.385 1.845 1.015 2.005 ;
        RECT  0.285 0.805 0.385 1.065 ;
        RECT  0.285 1.845 0.385 2.615 ;
        RECT  0.125 0.805 0.285 2.615 ;
    END
END DLY1X1

MACRO RFRDX4
    CLASS CORE ;
    FOREIGN RFRDX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.760 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 0.880 2.635 1.355 ;
        RECT  2.450 0.605 2.575 1.480 ;
        RECT  2.415 0.605 2.450 1.580 ;
        RECT  2.315 0.605 2.415 0.865 ;
        RECT  2.325 1.320 2.415 1.580 ;
        RECT  2.165 1.320 2.325 2.215 ;
        RECT  1.335 1.320 2.165 1.480 ;
        RECT  2.065 1.955 2.165 2.215 ;
        RECT  1.075 1.320 1.335 1.665 ;
        END
        ANTENNAGATEAREA     0.5512 ;
        ANTENNADIFFAREA     0.2715 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.625 1.660 1.885 2.050 ;
        RECT  0.900 1.850 1.625 2.050 ;
        RECT  0.895 0.540 0.900 1.140 ;
        RECT  0.895 1.850 0.900 2.895 ;
        RECT  0.640 0.540 0.895 2.895 ;
        RECT  0.585 0.695 0.640 2.585 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.8268 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 -0.250 2.760 0.250 ;
        RECT  1.185 -0.250 1.445 1.140 ;
        RECT  0.385 -0.250 1.185 0.250 ;
        RECT  0.125 -0.250 0.385 1.140 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 3.440 2.760 3.940 ;
        RECT  1.185 2.385 1.445 3.940 ;
        RECT  0.385 3.440 1.185 3.940 ;
        RECT  0.125 2.215 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
END RFRDX4

MACRO RFRDX2
    CLASS CORE ;
    FOREIGN RFRDX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 0.605 2.175 1.295 ;
        RECT  1.915 0.605 1.965 0.865 ;
        RECT  1.800 1.130 1.965 1.295 ;
        RECT  1.640 1.130 1.800 2.215 ;
        RECT  0.775 1.320 1.640 1.480 ;
        RECT  1.540 1.955 1.640 2.215 ;
        RECT  0.610 1.320 0.775 1.690 ;
        RECT  0.515 1.430 0.610 1.690 ;
        END
        ANTENNAGATEAREA     0.2756 ;
        ANTENNADIFFAREA     0.3208 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.100 1.660 1.360 2.030 ;
        RECT  0.385 1.870 1.100 2.030 ;
        RECT  0.335 0.625 0.385 1.225 ;
        RECT  0.335 1.870 0.385 3.045 ;
        RECT  0.125 0.625 0.335 3.045 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.7314 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 -0.250 2.300 0.250 ;
        RECT  0.670 -0.250 0.930 1.140 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 3.440 2.300 3.940 ;
        RECT  0.670 2.215 0.930 3.940 ;
        RECT  0.000 3.440 0.670 3.940 ;
        END
    END VDD
END RFRDX2

MACRO RFRDX1
    CLASS CORE ;
    FOREIGN RFRDX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.300 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 0.605 2.175 1.170 ;
        RECT  1.810 0.880 1.915 1.170 ;
        RECT  1.650 0.880 1.810 2.295 ;
        RECT  1.505 1.105 1.650 1.480 ;
        RECT  1.550 2.035 1.650 2.295 ;
        RECT  0.775 1.320 1.505 1.480 ;
        RECT  0.610 1.320 0.775 1.690 ;
        RECT  0.515 1.430 0.610 1.690 ;
        END
        ANTENNAGATEAREA     0.1378 ;
        ANTENNADIFFAREA     0.3209 ;
    END RB
    PIN BRB
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.110 1.665 1.370 2.035 ;
        RECT  0.385 1.875 1.110 2.035 ;
        RECT  0.335 0.990 0.385 1.250 ;
        RECT  0.335 1.875 0.385 2.555 ;
        RECT  0.125 0.990 0.335 2.555 ;
        END
        ANTENNAGATEAREA     0.1860 ;
        ANTENNADIFFAREA     0.3657 ;
    END BRB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 -0.250 2.300 0.250 ;
        RECT  0.670 -0.250 0.930 1.140 ;
        RECT  0.000 -0.250 0.670 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 3.440 2.300 3.940 ;
        RECT  0.670 2.215 0.930 3.940 ;
        RECT  0.000 3.440 0.670 3.940 ;
        END
    END VDD
END RFRDX1

MACRO RF2R1WX1
    CLASS CORE ;
    FOREIGN RF2R1WX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 2.930 2.635 3.220 ;
        RECT  2.325 2.930 2.425 3.150 ;
        RECT  2.065 2.890 2.325 3.150 ;
        END
        ANTENNAGATEAREA     0.1508 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.320 1.275 0.335 1.580 ;
        RECT  0.100 1.275 0.320 1.845 ;
        END
        ANTENNAGATEAREA     0.1807 ;
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.525 1.430 6.785 1.990 ;
        END
        ANTENNAGATEAREA     0.1716 ;
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 2.935 6.045 3.195 ;
        RECT  5.855 1.030 5.995 1.290 ;
        RECT  5.685 0.880 5.855 3.195 ;
        RECT  5.645 0.880 5.685 2.995 ;
        END
        ANTENNADIFFAREA     0.5490 ;
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.680 1.425 4.935 2.005 ;
        END
        ANTENNAGATEAREA     0.1742 ;
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.055 2.935 4.205 3.195 ;
        RECT  4.055 1.035 4.155 1.295 ;
        RECT  3.895 1.035 4.055 3.195 ;
        RECT  3.805 1.700 3.895 2.995 ;
        END
        ANTENNADIFFAREA     0.5536 ;
    END R1B
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.465 -0.250 6.900 0.250 ;
        RECT  6.205 -0.250 6.465 0.575 ;
        RECT  5.055 -0.250 6.205 0.250 ;
        RECT  4.795 -0.250 5.055 0.405 ;
        RECT  3.335 -0.250 4.795 0.250 ;
        RECT  3.175 -0.250 3.335 0.970 ;
        RECT  1.895 -0.250 3.175 0.250 ;
        RECT  1.635 -0.250 1.895 0.755 ;
        RECT  0.385 -0.250 1.635 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 3.440 6.900 3.940 ;
        RECT  6.305 2.895 6.565 3.940 ;
        RECT  5.000 3.440 6.305 3.940 ;
        RECT  5.000 2.860 5.170 3.120 ;
        RECT  4.740 2.860 5.000 3.940 ;
        RECT  4.570 2.860 4.740 3.120 ;
        RECT  3.370 3.440 4.740 3.940 ;
        RECT  3.110 2.390 3.370 3.940 ;
        RECT  1.885 3.440 3.110 3.940 ;
        RECT  1.625 2.690 1.885 3.940 ;
        RECT  0.385 3.440 1.625 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 1.025 6.565 1.185 ;
        RECT  6.345 2.265 6.565 2.525 ;
        RECT  6.305 1.025 6.345 2.525 ;
        RECT  6.185 1.025 6.305 2.475 ;
        RECT  6.180 1.745 6.185 2.475 ;
        RECT  6.045 1.745 6.180 2.005 ;
        RECT  5.275 1.400 5.395 1.660 ;
        RECT  5.115 0.685 5.275 1.660 ;
        RECT  3.715 0.685 5.115 0.845 ;
        RECT  4.495 1.085 4.715 1.245 ;
        RECT  4.455 2.275 4.715 2.535 ;
        RECT  4.400 1.085 4.495 1.650 ;
        RECT  4.415 2.275 4.455 2.435 ;
        RECT  4.400 1.905 4.415 2.435 ;
        RECT  4.335 1.085 4.400 2.435 ;
        RECT  4.240 1.490 4.335 2.435 ;
        RECT  3.555 0.685 3.715 1.435 ;
        RECT  3.530 1.275 3.555 1.435 ;
        RECT  3.410 1.275 3.530 1.760 ;
        RECT  3.250 1.275 3.410 2.180 ;
        RECT  2.855 1.275 3.250 1.435 ;
        RECT  2.860 2.020 3.250 2.180 ;
        RECT  2.070 1.615 3.015 1.775 ;
        RECT  2.700 2.020 2.860 2.750 ;
        RECT  2.595 1.035 2.855 1.435 ;
        RECT  2.600 2.490 2.700 2.750 ;
        RECT  1.730 1.275 2.595 1.435 ;
        RECT  2.240 0.525 2.475 0.785 ;
        RECT  2.250 1.955 2.410 2.510 ;
        RECT  1.440 2.350 2.250 2.510 ;
        RECT  2.215 0.525 2.240 1.095 ;
        RECT  2.080 0.575 2.215 1.095 ;
        RECT  1.390 0.935 2.080 1.095 ;
        RECT  1.910 1.615 2.070 2.170 ;
        RECT  1.100 2.010 1.910 2.170 ;
        RECT  1.570 1.275 1.730 1.830 ;
        RECT  1.280 2.350 1.440 3.040 ;
        RECT  1.230 0.695 1.390 1.095 ;
        RECT  0.925 2.880 1.280 3.040 ;
        RECT  0.675 0.695 1.230 0.855 ;
        RECT  1.050 2.010 1.100 2.700 ;
        RECT  0.890 1.035 1.050 2.700 ;
        RECT  0.665 2.880 0.925 3.140 ;
        RECT  0.840 2.100 0.890 2.700 ;
        RECT  0.660 0.695 0.675 1.920 ;
        RECT  0.660 2.880 0.665 3.040 ;
        RECT  0.515 0.695 0.660 3.040 ;
        RECT  0.500 1.760 0.515 3.040 ;
    END
END RF2R1WX1

MACRO RF1R1WX1
    CLASS CORE ;
    FOREIGN RF1R1WX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.680 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.520 1.715 2.810 ;
        RECT  1.260 2.550 1.505 2.810 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.370 1.580 0.400 1.840 ;
        RECT  0.125 1.505 0.370 1.990 ;
        END
        ANTENNAGATEAREA     0.0585 ;
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 2.110 3.555 2.555 ;
        RECT  3.245 2.140 3.275 2.400 ;
        END
        ANTENNAGATEAREA     0.0845 ;
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 0.945 3.200 1.305 ;
        RECT  2.885 0.880 3.095 1.305 ;
        END
        ANTENNAGATEAREA     0.0507 ;
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 2.735 3.555 2.995 ;
        RECT  3.380 0.505 3.540 1.930 ;
        RECT  3.275 0.505 3.380 0.765 ;
        RECT  3.060 1.770 3.380 1.930 ;
        RECT  3.060 2.735 3.295 2.895 ;
        RECT  2.900 1.770 3.060 2.895 ;
        RECT  2.425 2.520 2.900 2.810 ;
        END
        ANTENNADIFFAREA     0.3984 ;
    END RB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 -0.250 3.680 0.250 ;
        RECT  2.310 -0.250 2.570 0.795 ;
        RECT  0.390 -0.250 2.310 0.250 ;
        RECT  0.130 -0.250 0.390 0.795 ;
        RECT  0.000 -0.250 0.130 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 3.440 3.680 3.940 ;
        RECT  2.435 3.285 2.695 3.940 ;
        RECT  1.845 3.440 2.435 3.940 ;
        RECT  1.585 3.285 1.845 3.940 ;
        RECT  0.390 3.440 1.585 3.940 ;
        RECT  0.130 2.885 0.390 3.940 ;
        RECT  0.000 3.440 0.130 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.630 1.460 2.720 1.720 ;
        RECT  2.490 1.170 2.630 2.270 ;
        RECT  2.470 1.090 2.490 2.270 ;
        RECT  2.230 1.090 2.470 1.350 ;
        RECT  2.290 2.010 2.470 2.270 ;
        RECT  2.100 1.570 2.290 1.830 ;
        RECT  1.760 1.190 2.230 1.350 ;
        RECT  1.940 1.570 2.100 2.005 ;
        RECT  1.080 1.845 1.940 2.005 ;
        RECT  1.600 1.190 1.760 1.665 ;
        RECT  1.240 0.490 1.500 0.765 ;
        RECT  0.930 2.990 1.300 3.150 ;
        RECT  0.870 0.505 1.240 0.765 ;
        RECT  0.920 1.015 1.080 2.270 ;
        RECT  0.770 2.685 0.930 3.150 ;
        RECT  0.740 0.605 0.870 0.765 ;
        RECT  0.740 2.685 0.770 2.945 ;
        RECT  0.670 0.605 0.740 2.945 ;
        RECT  0.580 0.605 0.670 2.845 ;
    END
END RF1R1WX1

MACRO TLATNSRX4
    CLASS CORE ;
    FOREIGN TLATNSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.580 0.665 1.840 ;
        RECT  0.335 1.680 0.405 1.840 ;
        RECT  0.125 1.680 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 1.515 6.315 1.990 ;
        RECT  6.145 1.110 6.305 1.990 ;
        RECT  6.105 1.515 6.145 1.990 ;
        END
        ANTENNAGATEAREA     0.4186 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.865 1.105 10.915 2.400 ;
        RECT  10.605 0.655 10.865 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 1.700 9.995 2.400 ;
        RECT  9.585 0.655 9.845 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.885 1.370 7.145 1.630 ;
        RECT  6.775 1.370 6.885 1.580 ;
        RECT  6.565 1.290 6.775 1.580 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.455 4.545 1.615 ;
        RECT  2.475 1.455 2.635 1.990 ;
        RECT  2.425 1.545 2.475 1.990 ;
        RECT  2.350 1.545 2.425 1.805 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 -0.250 11.500 0.250 ;
        RECT  11.115 -0.250 11.375 1.190 ;
        RECT  10.355 -0.250 11.115 0.250 ;
        RECT  10.095 -0.250 10.355 1.205 ;
        RECT  9.305 -0.250 10.095 0.250 ;
        RECT  9.045 -0.250 9.305 0.405 ;
        RECT  8.535 -0.250 9.045 0.250 ;
        RECT  8.275 -0.250 8.535 0.405 ;
        RECT  7.045 -0.250 8.275 0.250 ;
        RECT  6.785 -0.250 7.045 0.405 ;
        RECT  4.345 -0.250 6.785 0.250 ;
        RECT  4.085 -0.250 4.345 0.590 ;
        RECT  1.005 -0.250 4.085 0.250 ;
        RECT  0.745 -0.250 1.005 0.815 ;
        RECT  0.000 -0.250 0.745 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.375 3.440 11.500 3.940 ;
        RECT  11.115 2.935 11.375 3.940 ;
        RECT  10.355 3.440 11.115 3.940 ;
        RECT  10.095 2.935 10.355 3.940 ;
        RECT  9.305 3.440 10.095 3.940 ;
        RECT  9.045 3.285 9.305 3.940 ;
        RECT  8.385 3.440 9.045 3.940 ;
        RECT  8.125 3.285 8.385 3.940 ;
        RECT  7.045 3.440 8.125 3.940 ;
        RECT  6.785 3.285 7.045 3.940 ;
        RECT  4.965 3.440 6.785 3.940 ;
        RECT  4.705 3.285 4.965 3.940 ;
        RECT  2.685 3.440 4.705 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  0.935 3.440 2.425 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.145 1.570 11.305 2.755 ;
        RECT  11.095 1.570 11.145 1.830 ;
        RECT  8.935 2.595 11.145 2.755 ;
        RECT  8.835 1.035 8.935 2.845 ;
        RECT  8.775 1.035 8.835 3.100 ;
        RECT  8.675 1.035 8.775 1.295 ;
        RECT  8.675 2.245 8.775 3.100 ;
        RECT  6.405 2.940 8.675 3.100 ;
        RECT  8.485 1.640 8.595 1.900 ;
        RECT  8.435 1.640 8.485 2.760 ;
        RECT  8.325 1.740 8.435 2.760 ;
        RECT  1.465 2.600 8.325 2.760 ;
        RECT  7.895 0.435 8.055 2.415 ;
        RECT  7.685 0.435 7.895 0.595 ;
        RECT  5.825 2.255 7.895 2.415 ;
        RECT  7.555 1.030 7.715 2.075 ;
        RECT  7.455 1.030 7.555 1.190 ;
        RECT  7.215 1.915 7.555 2.075 ;
        RECT  7.360 0.930 7.455 1.190 ;
        RECT  7.195 0.770 7.360 1.190 ;
        RECT  5.465 0.770 7.195 0.930 ;
        RECT  5.925 2.940 6.185 3.200 ;
        RECT  4.275 2.945 5.925 3.105 ;
        RECT  5.665 1.110 5.825 2.415 ;
        RECT  3.965 2.255 5.665 2.415 ;
        RECT  5.125 0.430 5.535 0.590 ;
        RECT  5.335 0.770 5.465 1.275 ;
        RECT  5.305 0.770 5.335 1.680 ;
        RECT  5.075 1.115 5.305 1.680 ;
        RECT  4.965 0.430 5.125 0.930 ;
        RECT  2.660 1.115 5.075 1.275 ;
        RECT  3.185 0.770 4.965 0.930 ;
        RECT  4.015 2.945 4.275 3.260 ;
        RECT  1.375 2.945 4.015 3.105 ;
        RECT  3.705 1.795 3.965 2.415 ;
        RECT  1.985 2.255 3.705 2.415 ;
        RECT  2.905 0.735 3.185 0.930 ;
        RECT  1.565 0.770 2.905 0.930 ;
        RECT  1.825 1.265 1.985 2.415 ;
        RECT  1.465 0.590 1.565 1.190 ;
        RECT  1.305 0.590 1.465 2.760 ;
        RECT  1.125 2.945 1.375 3.225 ;
        RECT  1.115 1.135 1.125 3.225 ;
        RECT  0.965 1.135 1.115 3.105 ;
        RECT  0.495 1.135 0.965 1.295 ;
        RECT  0.395 2.945 0.965 3.105 ;
        RECT  0.235 0.695 0.495 1.295 ;
        RECT  0.135 2.170 0.395 3.110 ;
    END
END TLATNSRX4

MACRO TLATNSRX2
    CLASS CORE ;
    FOREIGN TLATNSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.630 1.475 2.635 1.990 ;
        RECT  2.370 1.475 2.630 2.025 ;
        RECT  2.360 1.475 2.370 1.990 ;
        END
        ANTENNAGATEAREA     0.2288 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.655 7.695 3.060 ;
        RECT  7.435 0.655 7.535 1.255 ;
        RECT  7.435 2.120 7.535 3.060 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 1.515 6.775 2.400 ;
        RECT  6.565 1.035 6.615 2.400 ;
        RECT  6.465 1.035 6.565 2.335 ;
        RECT  6.455 1.035 6.465 2.215 ;
        RECT  6.355 1.035 6.455 1.295 ;
        RECT  6.415 1.955 6.455 2.215 ;
        END
        ANTENNADIFFAREA     0.6022 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.310 4.550 1.840 ;
        RECT  4.265 1.290 4.475 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.930 1.455 2.175 1.990 ;
        RECT  1.885 1.580 1.930 1.840 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 -0.250 7.820 0.250 ;
        RECT  6.895 -0.250 7.155 0.405 ;
        RECT  5.580 -0.250 6.895 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.500 -0.250 5.320 0.250 ;
        RECT  4.240 -0.250 4.500 0.405 ;
        RECT  2.065 -0.250 4.240 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 3.440 7.820 3.940 ;
        RECT  6.925 2.935 7.185 3.940 ;
        RECT  6.175 3.440 6.925 3.940 ;
        RECT  5.915 3.285 6.175 3.940 ;
        RECT  2.345 3.440 5.915 3.940 ;
        RECT  2.085 3.285 2.345 3.940 ;
        RECT  0.385 3.440 2.085 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.520 7.355 1.780 ;
        RECT  7.015 0.660 7.175 2.740 ;
        RECT  6.120 0.660 7.015 0.820 ;
        RECT  6.275 2.580 7.015 2.740 ;
        RECT  6.110 2.580 6.275 2.955 ;
        RECT  5.860 0.525 6.120 0.820 ;
        RECT  6.015 2.695 6.110 2.955 ;
        RECT  5.730 2.795 6.015 2.955 ;
        RECT  5.810 1.445 5.980 1.705 ;
        RECT  5.720 1.445 5.810 2.565 ;
        RECT  5.570 2.795 5.730 3.215 ;
        RECT  5.650 1.545 5.720 2.565 ;
        RECT  5.390 2.405 5.650 2.565 ;
        RECT  4.220 3.055 5.570 3.215 ;
        RECT  5.310 0.585 5.470 1.975 ;
        RECT  5.230 2.405 5.390 2.875 ;
        RECT  5.010 0.585 5.310 0.745 ;
        RECT  5.280 1.815 5.310 1.975 ;
        RECT  5.120 1.815 5.280 2.075 ;
        RECT  4.560 2.715 5.230 2.875 ;
        RECT  4.930 1.475 5.130 1.635 ;
        RECT  4.900 2.375 5.050 2.535 ;
        RECT  4.750 0.435 5.010 0.745 ;
        RECT  4.900 0.945 4.930 1.635 ;
        RECT  4.740 0.945 4.900 2.535 ;
        RECT  3.625 0.585 4.750 0.745 ;
        RECT  4.085 0.945 4.740 1.105 ;
        RECT  4.400 2.555 4.560 2.875 ;
        RECT  3.230 2.555 4.400 2.715 ;
        RECT  4.060 2.895 4.220 3.215 ;
        RECT  3.925 0.945 4.085 1.885 ;
        RECT  3.480 1.725 3.925 1.885 ;
        RECT  3.500 0.585 3.625 1.355 ;
        RECT  3.285 2.945 3.545 3.245 ;
        RECT  3.465 0.585 3.500 1.455 ;
        RECT  3.220 1.675 3.480 1.935 ;
        RECT  3.240 1.195 3.465 1.455 ;
        RECT  0.880 2.945 3.285 3.105 ;
        RECT  2.980 0.695 3.240 0.975 ;
        RECT  2.975 1.195 3.240 1.355 ;
        RECT  3.020 2.555 3.230 2.755 ;
        RECT  1.075 2.595 3.020 2.755 ;
        RECT  1.660 0.815 2.980 0.975 ;
        RECT  2.815 1.195 2.975 2.375 ;
        RECT  1.415 2.215 2.815 2.375 ;
        RECT  1.400 0.815 1.660 1.075 ;
        RECT  0.735 0.460 1.495 0.620 ;
        RECT  1.255 1.265 1.415 2.375 ;
        RECT  1.075 0.915 1.400 1.075 ;
        RECT  0.915 0.915 1.075 2.755 ;
        RECT  0.735 2.945 0.880 3.215 ;
        RECT  0.575 0.460 0.735 3.215 ;
    END
END TLATNSRX2

MACRO TLATNSRX1
    CLASS CORE ;
    FOREIGN TLATNSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.675 2.360 1.935 ;
        END
        ANTENNAGATEAREA     0.1391 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 0.880 6.775 2.330 ;
        RECT  6.615 0.845 6.655 2.330 ;
        RECT  6.565 0.845 6.615 1.170 ;
        RECT  6.565 1.925 6.615 2.330 ;
        RECT  6.395 0.845 6.565 1.105 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.3459 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.710 6.235 2.970 ;
        RECT  5.870 2.710 5.975 2.870 ;
        RECT  5.710 1.035 5.870 2.870 ;
        END
        ANTENNADIFFAREA     0.3276 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.470 4.325 1.730 ;
        RECT  3.825 1.470 4.015 1.990 ;
        RECT  3.805 1.700 3.825 1.990 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.600 2.005 1.860 ;
        RECT  1.745 1.420 1.905 1.860 ;
        RECT  1.715 1.420 1.745 1.580 ;
        RECT  1.505 1.290 1.715 1.580 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.080 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.385 3.440 4.220 3.940 ;
        RECT  2.125 3.285 2.385 3.940 ;
        RECT  0.385 3.440 2.125 3.940 ;
        RECT  0.125 2.870 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.210 1.360 6.435 1.520 ;
        RECT  6.050 0.590 6.210 1.520 ;
        RECT  5.890 0.590 6.050 0.750 ;
        RECT  5.630 0.465 5.890 0.750 ;
        RECT  5.490 0.590 5.630 0.750 ;
        RECT  5.490 1.600 5.530 2.900 ;
        RECT  5.370 0.590 5.490 2.900 ;
        RECT  5.330 0.590 5.370 1.760 ;
        RECT  4.990 2.740 5.370 2.900 ;
        RECT  5.145 1.955 5.190 2.215 ;
        RECT  4.985 0.690 5.145 2.215 ;
        RECT  4.300 2.400 5.040 2.560 ;
        RECT  4.725 2.740 4.990 3.105 ;
        RECT  4.725 0.690 4.985 0.850 ;
        RECT  4.705 1.080 4.805 2.215 ;
        RECT  4.465 0.490 4.725 0.850 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.645 1.030 4.705 2.215 ;
        RECT  4.445 1.030 4.645 1.290 ;
        RECT  4.470 1.955 4.645 2.215 ;
        RECT  3.285 0.690 4.465 0.850 ;
        RECT  3.625 1.130 4.445 1.290 ;
        RECT  4.140 2.400 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.485 1.130 3.625 2.000 ;
        RECT  3.465 1.130 3.485 2.100 ;
        RECT  3.225 1.840 3.465 2.100 ;
        RECT  3.125 0.690 3.285 1.625 ;
        RECT  3.015 1.410 3.125 1.625 ;
        RECT  2.975 1.465 3.015 1.625 ;
        RECT  2.815 1.465 2.975 2.335 ;
        RECT  2.785 0.950 2.945 1.225 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.475 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.785 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  1.215 0.510 1.475 0.770 ;
        RECT  1.315 1.760 1.475 2.335 ;
        RECT  1.105 0.950 1.325 1.270 ;
        RECT  0.765 0.610 1.215 0.770 ;
        RECT  1.105 2.535 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.575 2.745 0.605 3.005 ;
    END
END TLATNSRX1

MACRO TLATNSRXL
    CLASS CORE ;
    FOREIGN TLATNSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.850 ;
        RECT  0.125 1.290 0.335 1.850 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.765 2.360 1.925 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.175 ;
        RECT  6.565 0.865 6.725 2.330 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.2585 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.730 6.235 3.010 ;
        RECT  5.870 1.020 6.030 1.280 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.020 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.470 4.375 1.730 ;
        RECT  3.805 1.290 4.015 1.730 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.290 2.175 1.580 ;
        RECT  1.925 1.420 1.965 1.580 ;
        RECT  1.765 1.420 1.925 1.965 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.070 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.235 3.440 4.220 3.940 ;
        RECT  1.975 3.285 2.235 3.940 ;
        RECT  0.385 3.440 1.975 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 0.610 6.385 1.495 ;
        RECT  6.030 0.610 6.225 0.770 ;
        RECT  5.770 0.510 6.030 0.770 ;
        RECT  5.530 0.610 5.770 0.770 ;
        RECT  5.370 0.610 5.530 2.890 ;
        RECT  4.990 2.730 5.370 2.890 ;
        RECT  5.030 0.690 5.190 2.215 ;
        RECT  4.725 0.690 5.030 0.850 ;
        RECT  4.725 2.730 4.990 3.105 ;
        RECT  4.300 2.390 4.850 2.550 ;
        RECT  4.645 1.030 4.805 2.165 ;
        RECT  4.465 0.520 4.725 0.850 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.445 1.030 4.645 1.290 ;
        RECT  3.415 2.005 4.645 2.165 ;
        RECT  3.505 0.690 4.465 0.850 ;
        RECT  4.140 2.390 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.345 0.690 3.505 1.570 ;
        RECT  3.155 1.840 3.415 2.165 ;
        RECT  2.975 1.410 3.345 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.335 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.445 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  0.765 0.610 1.535 0.770 ;
        RECT  1.285 1.705 1.445 2.335 ;
        RECT  1.105 0.950 1.325 1.250 ;
        RECT  1.105 2.535 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.600 2.685 0.605 2.945 ;
    END
END TLATNSRXL

MACRO TLATNX4
    CLASS CORE ;
    FOREIGN TLATNX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 1.105 6.775 1.990 ;
        RECT  6.465 0.695 6.725 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 1.290 5.855 1.990 ;
        RECT  5.445 0.695 5.705 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.895 ;
        RECT  0.110 1.515 0.125 1.895 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.485 1.835 1.990 ;
        RECT  1.505 1.700 1.575 1.990 ;
        END
        ANTENNAGATEAREA     0.4628 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 -0.250 7.360 0.250 ;
        RECT  6.975 -0.250 7.235 1.095 ;
        RECT  6.215 -0.250 6.975 0.250 ;
        RECT  5.955 -0.250 6.215 1.095 ;
        RECT  5.190 -0.250 5.955 0.250 ;
        RECT  4.930 -0.250 5.190 1.095 ;
        RECT  3.485 -0.250 4.930 0.250 ;
        RECT  3.225 -0.250 3.485 0.405 ;
        RECT  1.695 -0.250 3.225 0.250 ;
        RECT  1.435 -0.250 1.695 0.735 ;
        RECT  0.385 -0.250 1.435 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 3.440 7.360 3.940 ;
        RECT  6.975 2.940 7.235 3.940 ;
        RECT  6.215 3.440 6.975 3.940 ;
        RECT  5.955 2.940 6.215 3.940 ;
        RECT  5.165 3.440 5.955 3.940 ;
        RECT  4.905 3.285 5.165 3.940 ;
        RECT  3.220 3.440 4.905 3.940 ;
        RECT  3.060 2.955 3.220 3.940 ;
        RECT  1.580 3.440 3.060 3.940 ;
        RECT  1.320 2.955 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.150 1.580 7.250 1.840 ;
        RECT  6.990 1.580 7.150 2.760 ;
        RECT  5.225 2.600 6.990 2.760 ;
        RECT  5.065 1.280 5.225 2.760 ;
        RECT  4.725 1.280 5.065 1.440 ;
        RECT  4.725 2.600 5.065 2.760 ;
        RECT  4.355 1.795 4.885 2.055 ;
        RECT  4.610 0.655 4.725 1.440 ;
        RECT  4.465 2.600 4.725 2.910 ;
        RECT  4.565 0.555 4.610 1.440 ;
        RECT  4.350 0.555 4.565 0.815 ;
        RECT  3.590 2.750 4.465 2.910 ;
        RECT  4.270 1.115 4.355 2.055 ;
        RECT  3.985 0.655 4.350 0.815 ;
        RECT  4.195 1.115 4.270 2.420 ;
        RECT  3.475 1.115 4.195 1.275 ;
        RECT  4.110 1.895 4.195 2.420 ;
        RECT  3.175 2.260 4.110 2.420 ;
        RECT  3.855 1.455 4.015 1.715 ;
        RECT  3.725 0.475 3.985 0.815 ;
        RECT  3.135 1.455 3.855 1.615 ;
        RECT  3.430 2.750 3.590 3.120 ;
        RECT  2.795 1.815 3.585 1.975 ;
        RECT  3.315 0.795 3.475 1.275 ;
        RECT  2.585 0.795 3.315 0.955 ;
        RECT  3.015 2.260 3.175 2.775 ;
        RECT  2.975 1.145 3.135 1.615 ;
        RECT  2.435 2.615 3.015 2.775 ;
        RECT  2.215 1.145 2.975 1.305 ;
        RECT  2.695 1.485 2.795 1.975 ;
        RECT  2.535 1.485 2.695 2.410 ;
        RECT  2.325 0.695 2.585 0.955 ;
        RECT  1.995 2.250 2.535 2.410 ;
        RECT  2.175 2.615 2.435 3.215 ;
        RECT  2.215 1.805 2.315 2.065 ;
        RECT  2.055 1.145 2.215 2.065 ;
        RECT  1.265 1.145 2.055 1.305 ;
        RECT  1.835 2.250 1.995 2.740 ;
        RECT  0.785 2.580 1.835 2.740 ;
        RECT  1.185 1.140 1.265 2.400 ;
        RECT  1.105 0.525 1.185 2.400 ;
        RECT  1.025 0.525 1.105 1.305 ;
        RECT  0.925 2.140 1.105 2.400 ;
        RECT  0.925 0.525 1.025 0.785 ;
        RECT  0.710 1.640 0.925 1.900 ;
        RECT  0.710 1.035 0.815 1.295 ;
        RECT  0.710 2.580 0.785 2.910 ;
        RECT  0.550 1.035 0.710 2.910 ;
        RECT  0.525 2.650 0.550 2.910 ;
    END
END TLATNX4

MACRO TLATNX2
    CLASS CORE ;
    FOREIGN TLATNX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.390 0.695 5.395 0.945 ;
        RECT  5.390 2.335 5.395 2.995 ;
        RECT  5.230 0.575 5.390 3.045 ;
        RECT  5.130 0.575 5.230 1.175 ;
        RECT  5.130 2.105 5.230 3.045 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.515 4.475 1.990 ;
        RECT  4.310 1.515 4.340 2.900 ;
        RECT  4.080 1.035 4.310 2.900 ;
        RECT  4.050 1.035 4.080 1.295 ;
        END
        ANTENNADIFFAREA     0.6988 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.335 1.260 0.360 1.735 ;
        RECT  0.125 1.260 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0832 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 1.290 1.715 1.580 ;
        RECT  1.395 1.085 1.680 1.600 ;
        END
        ANTENNAGATEAREA     0.2522 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 -0.250 5.520 0.250 ;
        RECT  4.590 -0.250 4.850 0.405 ;
        RECT  3.260 -0.250 4.590 0.250 ;
        RECT  3.000 -0.250 3.260 0.925 ;
        RECT  1.465 -0.250 3.000 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.850 3.440 5.520 3.940 ;
        RECT  4.590 2.245 4.850 3.940 ;
        RECT  3.220 3.440 4.590 3.940 ;
        RECT  2.960 2.485 3.220 3.940 ;
        RECT  1.360 3.440 2.960 3.940 ;
        RECT  1.100 3.285 1.360 3.940 ;
        RECT  0.385 3.440 1.100 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.950 1.405 5.050 1.665 ;
        RECT  4.790 0.695 4.950 1.665 ;
        RECT  3.800 0.695 4.790 0.855 ;
        RECT  3.705 2.420 3.830 2.680 ;
        RECT  3.705 0.695 3.800 1.005 ;
        RECT  3.545 0.695 3.705 2.680 ;
        RECT  3.540 0.695 3.545 1.005 ;
        RECT  2.960 1.990 3.545 2.250 ;
        RECT  2.780 1.220 3.365 1.480 ;
        RECT  2.620 1.220 2.780 2.755 ;
        RECT  2.315 1.220 2.620 1.380 ;
        RECT  2.230 2.595 2.620 2.755 ;
        RECT  2.315 0.445 2.575 0.745 ;
        RECT  2.280 2.145 2.440 2.410 ;
        RECT  1.215 0.585 2.315 0.745 ;
        RECT  2.155 0.965 2.315 1.380 ;
        RECT  1.715 2.250 2.280 2.410 ;
        RECT  1.970 2.595 2.230 3.195 ;
        RECT  2.055 0.965 2.155 1.225 ;
        RECT  1.895 1.665 2.155 1.945 ;
        RECT  1.215 1.785 1.895 1.945 ;
        RECT  1.555 2.250 1.715 3.105 ;
        RECT  0.380 2.945 1.555 3.105 ;
        RECT  1.055 0.585 1.215 2.765 ;
        RECT  0.895 0.585 1.055 0.785 ;
        RECT  0.560 2.605 1.055 2.765 ;
        RECT  0.635 0.525 0.895 0.785 ;
        RECT  0.815 1.515 0.875 1.840 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.525 1.955 0.655 2.330 ;
        RECT  0.380 2.170 0.525 2.330 ;
        RECT  0.220 2.170 0.380 3.105 ;
    END
END TLATNX2

MACRO TLATNX1
    CLASS CORE ;
    FOREIGN TLATNX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.025 4.475 2.810 ;
        RECT  4.255 1.025 4.265 1.285 ;
        RECT  4.215 2.305 4.265 2.565 ;
        END
        ANTENNADIFFAREA     0.4535 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.035 0.595 4.075 2.125 ;
        RECT  3.915 0.595 4.035 2.855 ;
        RECT  3.680 0.595 3.915 0.755 ;
        RECT  3.875 1.965 3.915 2.855 ;
        RECT  3.805 2.520 3.875 2.855 ;
        RECT  3.250 2.595 3.805 2.855 ;
        RECT  3.420 0.430 3.680 0.755 ;
        END
        ANTENNADIFFAREA     0.3691 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.335 1.260 0.360 1.735 ;
        RECT  0.125 1.260 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 1.290 1.715 1.580 ;
        RECT  1.395 1.080 1.680 1.595 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 -0.250 4.600 0.250 ;
        RECT  4.010 -0.250 4.270 0.405 ;
        RECT  3.055 -0.250 4.010 0.250 ;
        RECT  2.795 -0.250 3.055 0.405 ;
        RECT  1.475 -0.250 2.795 0.250 ;
        RECT  1.215 -0.250 1.475 0.405 ;
        RECT  0.385 -0.250 1.215 0.250 ;
        RECT  0.125 -0.250 0.385 0.805 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 3.440 4.600 3.940 ;
        RECT  3.620 3.285 3.880 3.940 ;
        RECT  2.925 3.440 3.620 3.940 ;
        RECT  2.665 3.285 2.925 3.940 ;
        RECT  1.325 3.440 2.665 3.940 ;
        RECT  1.065 3.065 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.635 1.500 3.735 1.760 ;
        RECT  3.475 1.125 3.635 2.295 ;
        RECT  3.375 1.125 3.475 1.385 ;
        RECT  2.985 2.135 3.475 2.295 ;
        RECT  2.645 1.685 3.255 1.945 ;
        RECT  2.825 2.135 2.985 3.075 ;
        RECT  2.375 2.915 2.825 3.075 ;
        RECT  2.485 1.025 2.645 2.435 ;
        RECT  2.255 0.485 2.515 0.745 ;
        RECT  2.285 1.025 2.485 1.185 ;
        RECT  2.065 2.275 2.485 2.435 ;
        RECT  2.025 0.925 2.285 1.185 ;
        RECT  1.215 0.585 2.255 0.745 ;
        RECT  1.805 2.175 2.065 2.435 ;
        RECT  1.215 1.775 1.905 1.935 ;
        RECT  1.055 0.585 1.215 2.555 ;
        RECT  0.895 0.585 1.055 0.785 ;
        RECT  0.745 2.395 1.055 2.555 ;
        RECT  0.635 0.525 0.895 0.785 ;
        RECT  0.815 1.515 0.875 1.840 ;
        RECT  0.655 1.035 0.815 2.215 ;
        RECT  0.585 2.395 0.745 2.815 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.525 1.955 0.655 2.215 ;
        RECT  0.485 2.555 0.585 2.815 ;
    END
END TLATNX1

MACRO TLATNXL
    CLASS CORE ;
    FOREIGN TLATNXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.265 1.025 4.475 2.565 ;
        RECT  4.215 2.305 4.265 2.565 ;
        END
        ANTENNADIFFAREA     0.2827 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 0.625 4.075 2.125 ;
        RECT  3.915 0.625 3.970 2.680 ;
        RECT  3.680 0.625 3.915 0.785 ;
        RECT  3.810 1.965 3.915 2.680 ;
        RECT  3.555 2.520 3.810 2.680 ;
        RECT  3.420 0.525 3.680 0.785 ;
        RECT  3.510 2.520 3.555 2.810 ;
        RECT  3.250 2.520 3.510 2.855 ;
        END
        ANTENNADIFFAREA     0.2340 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.475 0.445 1.735 ;
        RECT  0.125 1.300 0.360 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.670 1.290 1.715 1.580 ;
        RECT  1.395 1.080 1.670 1.595 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 -0.250 4.600 0.250 ;
        RECT  4.020 -0.250 4.280 0.405 ;
        RECT  3.095 -0.250 4.020 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  1.465 -0.250 2.835 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.805 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 3.440 4.600 3.940 ;
        RECT  3.620 3.285 3.880 3.940 ;
        RECT  3.035 3.440 3.620 3.940 ;
        RECT  2.775 3.285 3.035 3.940 ;
        RECT  1.385 3.440 2.775 3.940 ;
        RECT  1.125 3.285 1.385 3.940 ;
        RECT  0.385 3.440 1.125 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.630 1.500 3.735 1.760 ;
        RECT  3.630 1.035 3.680 1.295 ;
        RECT  3.470 1.035 3.630 2.295 ;
        RECT  3.420 1.035 3.470 1.295 ;
        RECT  2.985 2.135 3.470 2.295 ;
        RECT  2.870 1.685 3.255 1.945 ;
        RECT  2.825 2.135 2.985 3.060 ;
        RECT  2.710 0.735 2.870 1.945 ;
        RECT  2.595 2.900 2.825 3.060 ;
        RECT  2.315 0.735 2.710 0.895 ;
        RECT  2.645 1.785 2.710 1.945 ;
        RECT  2.485 1.785 2.645 2.370 ;
        RECT  2.335 2.900 2.595 3.160 ;
        RECT  2.305 1.080 2.515 1.240 ;
        RECT  2.125 2.210 2.485 2.370 ;
        RECT  2.055 0.635 2.315 0.895 ;
        RECT  2.145 1.080 2.305 2.030 ;
        RECT  1.215 1.870 2.145 2.030 ;
        RECT  1.865 2.210 2.125 2.470 ;
        RECT  1.810 2.900 2.070 3.160 ;
        RECT  0.305 2.945 1.810 3.105 ;
        RECT  1.055 0.590 1.215 2.765 ;
        RECT  0.895 0.590 1.055 0.750 ;
        RECT  0.485 2.605 1.055 2.765 ;
        RECT  0.635 0.430 0.895 0.750 ;
        RECT  0.815 1.515 0.875 1.780 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.555 1.960 0.655 2.330 ;
        RECT  0.305 2.170 0.555 2.330 ;
        RECT  0.145 2.170 0.305 3.105 ;
    END
END TLATNXL

MACRO TLATSRX4
    CLASS CORE ;
    FOREIGN TLATSRX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.500 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.580 0.665 1.860 ;
        RECT  0.335 1.700 0.405 1.860 ;
        RECT  0.125 1.700 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.2561 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.195 6.405 1.730 ;
        END
        ANTENNAGATEAREA     0.4212 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.855 1.105 10.915 2.400 ;
        RECT  10.595 0.655 10.855 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.835 1.700 9.995 2.400 ;
        RECT  9.575 0.655 9.835 2.400 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.855 1.290 7.235 1.665 ;
        END
        ANTENNAGATEAREA     0.1443 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.445 1.445 4.705 1.615 ;
        RECT  2.745 1.445 4.445 1.605 ;
        RECT  2.635 1.445 2.745 1.925 ;
        RECT  2.585 1.445 2.635 1.990 ;
        RECT  2.485 1.535 2.585 1.990 ;
        RECT  2.425 1.700 2.485 1.990 ;
        END
        ANTENNAGATEAREA     0.4264 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.365 -0.250 11.500 0.250 ;
        RECT  11.105 -0.250 11.365 1.190 ;
        RECT  10.345 -0.250 11.105 0.250 ;
        RECT  10.085 -0.250 10.345 1.205 ;
        RECT  9.285 -0.250 10.085 0.250 ;
        RECT  9.025 -0.250 9.285 0.405 ;
        RECT  8.525 -0.250 9.025 0.250 ;
        RECT  8.265 -0.250 8.525 0.405 ;
        RECT  7.145 -0.250 8.265 0.250 ;
        RECT  6.885 -0.250 7.145 0.405 ;
        RECT  4.500 -0.250 6.885 0.250 ;
        RECT  4.240 -0.250 4.500 0.585 ;
        RECT  0.935 -0.250 4.240 0.250 ;
        RECT  0.675 -0.250 0.935 0.945 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.370 3.440 11.500 3.940 ;
        RECT  11.110 2.935 11.370 3.940 ;
        RECT  10.345 3.440 11.110 3.940 ;
        RECT  10.085 2.935 10.345 3.940 ;
        RECT  9.285 3.440 10.085 3.940 ;
        RECT  9.025 3.285 9.285 3.940 ;
        RECT  8.365 3.440 9.025 3.940 ;
        RECT  8.105 3.285 8.365 3.940 ;
        RECT  7.040 3.440 8.105 3.940 ;
        RECT  6.780 3.285 7.040 3.940 ;
        RECT  4.815 3.440 6.780 3.940 ;
        RECT  4.555 3.285 4.815 3.940 ;
        RECT  2.685 3.440 4.555 3.940 ;
        RECT  2.425 3.285 2.685 3.940 ;
        RECT  0.935 3.440 2.425 3.940 ;
        RECT  0.675 3.285 0.935 3.940 ;
        RECT  0.000 3.440 0.675 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.095 1.570 11.255 2.755 ;
        RECT  8.925 2.595 11.095 2.755 ;
        RECT  8.825 1.035 8.925 2.845 ;
        RECT  8.765 1.035 8.825 3.105 ;
        RECT  8.665 1.035 8.765 1.295 ;
        RECT  8.665 2.245 8.765 3.105 ;
        RECT  6.410 2.945 8.665 3.105 ;
        RECT  8.485 1.785 8.585 2.045 ;
        RECT  8.325 1.785 8.485 2.760 ;
        RECT  1.520 2.600 8.325 2.760 ;
        RECT  7.935 0.610 8.085 2.370 ;
        RECT  7.925 0.435 7.935 2.370 ;
        RECT  7.675 0.435 7.925 0.770 ;
        RECT  7.690 2.210 7.925 2.370 ;
        RECT  7.575 1.470 7.745 1.730 ;
        RECT  7.000 0.610 7.675 0.770 ;
        RECT  7.440 0.950 7.575 2.005 ;
        RECT  7.415 0.950 7.440 2.415 ;
        RECT  7.285 0.950 7.415 1.110 ;
        RECT  7.280 1.845 7.415 2.415 ;
        RECT  7.180 2.115 7.280 2.415 ;
        RECT  5.925 2.255 7.180 2.415 ;
        RECT  6.840 0.610 7.000 0.935 ;
        RECT  5.575 0.775 6.840 0.935 ;
        RECT  4.275 2.945 6.190 3.105 ;
        RECT  5.765 1.115 5.925 2.415 ;
        RECT  3.965 2.255 5.765 2.415 ;
        RECT  5.235 0.430 5.705 0.590 ;
        RECT  5.495 0.775 5.575 1.265 ;
        RECT  5.415 0.775 5.495 1.685 ;
        RECT  5.235 1.105 5.415 1.685 ;
        RECT  5.075 0.430 5.235 0.925 ;
        RECT  3.055 1.105 5.235 1.265 ;
        RECT  3.440 0.765 5.075 0.925 ;
        RECT  4.015 2.945 4.275 3.235 ;
        RECT  1.375 2.945 4.015 3.105 ;
        RECT  3.705 1.785 3.965 2.415 ;
        RECT  2.105 2.255 3.705 2.415 ;
        RECT  3.280 0.665 3.440 0.925 ;
        RECT  1.520 0.665 3.280 0.825 ;
        RECT  2.795 1.005 3.055 1.265 ;
        RECT  1.945 1.250 2.105 2.415 ;
        RECT  1.360 0.625 1.520 2.760 ;
        RECT  1.115 2.945 1.375 3.230 ;
        RECT  1.185 0.625 1.360 1.225 ;
        RECT  1.255 2.160 1.360 2.760 ;
        RECT  1.005 1.405 1.180 1.665 ;
        RECT  1.005 2.945 1.115 3.105 ;
        RECT  0.845 1.135 1.005 3.105 ;
        RECT  0.425 1.135 0.845 1.295 ;
        RECT  0.385 2.945 0.845 3.105 ;
        RECT  0.165 0.695 0.425 1.295 ;
        RECT  0.125 2.170 0.385 3.110 ;
    END
END TLATSRX4

MACRO TLATSRX2
    CLASS CORE ;
    FOREIGN TLATSRX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.820 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 2.025 ;
        END
        ANTENNAGATEAREA     0.2288 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 0.655 7.695 3.060 ;
        RECT  7.435 0.655 7.535 1.255 ;
        RECT  7.435 2.120 7.535 3.060 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 1.515 6.775 2.400 ;
        RECT  6.565 1.035 6.615 2.400 ;
        RECT  6.455 1.035 6.565 2.215 ;
        RECT  6.355 1.035 6.455 1.295 ;
        RECT  6.415 1.955 6.455 2.215 ;
        END
        ANTENNADIFFAREA     0.5833 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.475 1.310 4.550 1.840 ;
        RECT  4.265 1.290 4.475 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.290 2.175 1.845 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 -0.250 7.820 0.250 ;
        RECT  6.895 -0.250 7.155 0.405 ;
        RECT  5.580 -0.250 6.895 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.500 -0.250 5.320 0.250 ;
        RECT  4.240 -0.250 4.500 0.405 ;
        RECT  2.065 -0.250 4.240 0.250 ;
        RECT  1.805 -0.250 2.065 0.405 ;
        RECT  0.385 -0.250 1.805 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 3.440 7.820 3.940 ;
        RECT  6.925 2.935 7.185 3.940 ;
        RECT  6.175 3.440 6.925 3.940 ;
        RECT  5.915 3.285 6.175 3.940 ;
        RECT  2.345 3.440 5.915 3.940 ;
        RECT  2.085 3.285 2.345 3.940 ;
        RECT  0.385 3.440 2.085 3.940 ;
        RECT  0.125 2.945 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.175 1.520 7.355 1.780 ;
        RECT  7.015 0.660 7.175 2.740 ;
        RECT  6.150 0.660 7.015 0.820 ;
        RECT  6.275 2.580 7.015 2.740 ;
        RECT  6.175 2.465 6.275 2.740 ;
        RECT  6.015 2.465 6.175 2.955 ;
        RECT  5.890 0.525 6.150 0.820 ;
        RECT  5.730 2.795 6.015 2.955 ;
        RECT  5.810 1.445 5.980 1.705 ;
        RECT  5.720 1.445 5.810 2.565 ;
        RECT  5.570 2.795 5.730 3.215 ;
        RECT  5.650 1.545 5.720 2.565 ;
        RECT  5.390 2.405 5.650 2.565 ;
        RECT  4.220 3.055 5.570 3.215 ;
        RECT  5.310 0.865 5.470 1.975 ;
        RECT  5.230 2.405 5.390 2.875 ;
        RECT  5.295 0.865 5.310 1.025 ;
        RECT  5.280 1.815 5.310 1.975 ;
        RECT  5.135 0.585 5.295 1.025 ;
        RECT  5.120 1.815 5.280 2.075 ;
        RECT  4.560 2.715 5.230 2.875 ;
        RECT  5.010 0.585 5.135 0.745 ;
        RECT  4.930 1.475 5.130 1.635 ;
        RECT  4.900 2.375 5.050 2.535 ;
        RECT  4.750 0.435 5.010 0.745 ;
        RECT  4.900 0.945 4.930 1.635 ;
        RECT  4.740 0.945 4.900 2.535 ;
        RECT  4.085 0.585 4.750 0.745 ;
        RECT  4.670 0.945 4.740 1.105 ;
        RECT  2.975 2.215 4.740 2.375 ;
        RECT  4.400 2.555 4.560 2.875 ;
        RECT  1.075 2.555 4.400 2.715 ;
        RECT  4.060 2.895 4.220 3.215 ;
        RECT  3.925 0.585 4.085 1.835 ;
        RECT  3.480 1.675 3.925 1.835 ;
        RECT  3.285 2.945 3.545 3.245 ;
        RECT  2.975 1.195 3.500 1.455 ;
        RECT  3.220 1.675 3.480 1.935 ;
        RECT  0.880 2.945 3.285 3.105 ;
        RECT  2.980 0.695 3.240 0.975 ;
        RECT  1.660 0.815 2.980 0.975 ;
        RECT  2.815 1.195 2.975 2.375 ;
        RECT  1.415 2.215 2.815 2.375 ;
        RECT  1.400 0.815 1.660 1.075 ;
        RECT  0.735 0.460 1.495 0.620 ;
        RECT  1.255 1.265 1.415 2.375 ;
        RECT  1.075 0.915 1.400 1.075 ;
        RECT  0.915 0.915 1.075 2.715 ;
        RECT  0.735 2.945 0.880 3.255 ;
        RECT  0.575 0.460 0.735 3.255 ;
    END
END TLATSRX2

MACRO TLATSRX1
    CLASS CORE ;
    FOREIGN TLATSRX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.840 ;
        RECT  0.125 1.290 0.335 1.840 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.675 2.360 1.935 ;
        END
        ANTENNAGATEAREA     0.1391 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.180 ;
        RECT  6.565 0.880 6.725 2.330 ;
        RECT  6.395 0.895 6.565 1.055 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.3459 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  6.135 2.950 6.235 3.210 ;
        RECT  5.975 2.730 6.135 3.210 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.035 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.3276 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 1.420 4.325 1.705 ;
        RECT  4.015 1.375 4.260 1.705 ;
        RECT  3.805 1.290 4.015 1.705 ;
        END
        ANTENNAGATEAREA     0.0689 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 1.600 2.005 1.860 ;
        RECT  1.745 1.420 1.905 1.860 ;
        RECT  1.715 1.420 1.745 1.580 ;
        RECT  1.505 1.290 1.715 1.580 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.695 3.440 6.515 3.940 ;
        RECT  5.435 3.080 5.695 3.940 ;
        RECT  4.470 3.440 5.435 3.940 ;
        RECT  4.210 3.285 4.470 3.940 ;
        RECT  2.380 3.440 4.210 3.940 ;
        RECT  2.120 3.285 2.380 3.940 ;
        RECT  0.385 3.440 2.120 3.940 ;
        RECT  0.125 2.870 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 1.260 6.385 1.520 ;
        RECT  6.210 1.260 6.225 1.420 ;
        RECT  6.050 0.590 6.210 1.420 ;
        RECT  5.890 0.590 6.050 0.750 ;
        RECT  5.630 0.465 5.890 0.750 ;
        RECT  5.490 0.590 5.630 0.750 ;
        RECT  5.490 1.600 5.530 2.900 ;
        RECT  5.370 0.590 5.490 2.900 ;
        RECT  5.330 0.590 5.370 1.760 ;
        RECT  5.120 2.740 5.370 2.900 ;
        RECT  5.145 1.955 5.190 2.215 ;
        RECT  4.985 0.700 5.145 2.215 ;
        RECT  4.860 2.740 5.120 3.105 ;
        RECT  4.300 2.400 5.040 2.560 ;
        RECT  4.725 0.700 4.985 0.860 ;
        RECT  4.030 2.945 4.860 3.105 ;
        RECT  4.645 1.080 4.805 2.215 ;
        RECT  4.465 0.520 4.725 0.860 ;
        RECT  4.445 1.080 4.645 1.240 ;
        RECT  4.470 1.955 4.645 2.215 ;
        RECT  3.960 2.055 4.470 2.215 ;
        RECT  3.615 0.700 4.465 0.860 ;
        RECT  4.140 2.400 4.300 2.745 ;
        RECT  1.210 2.585 4.140 2.745 ;
        RECT  3.870 2.945 4.030 3.255 ;
        RECT  3.800 2.055 3.960 2.405 ;
        RECT  2.975 2.245 3.800 2.405 ;
        RECT  3.455 0.700 3.615 2.050 ;
        RECT  3.155 1.890 3.455 2.050 ;
        RECT  2.975 1.410 3.275 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.405 ;
        RECT  2.660 2.945 2.920 3.255 ;
        RECT  1.475 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.755 2.945 2.660 3.105 ;
        RECT  1.215 0.510 1.475 0.770 ;
        RECT  1.315 1.760 1.475 2.335 ;
        RECT  1.105 0.950 1.325 1.270 ;
        RECT  0.740 0.610 1.215 0.770 ;
        RECT  1.105 2.515 1.210 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.740 1.035 0.765 1.295 ;
        RECT  0.740 2.795 0.755 3.105 ;
        RECT  0.595 0.610 0.740 3.105 ;
        RECT  0.580 0.610 0.595 3.005 ;
        RECT  0.565 2.745 0.580 3.005 ;
    END
END TLATSRX1

MACRO TLATSRXL
    CLASS CORE ;
    FOREIGN TLATSRXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.900 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.355 0.395 1.850 ;
        RECT  0.125 1.290 0.335 1.850 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.475 2.635 1.990 ;
        RECT  2.225 1.760 2.360 1.920 ;
        END
        ANTENNAGATEAREA     0.1014 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.725 0.880 6.775 2.175 ;
        RECT  6.565 0.865 6.725 2.330 ;
        RECT  6.215 2.170 6.565 2.330 ;
        RECT  6.055 2.170 6.215 2.430 ;
        END
        ANTENNADIFFAREA     0.2585 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.870 1.700 6.315 1.990 ;
        RECT  5.975 2.730 6.235 3.010 ;
        RECT  5.870 1.020 6.030 1.280 ;
        RECT  5.870 2.730 5.975 2.890 ;
        RECT  5.710 1.020 5.870 2.890 ;
        END
        ANTENNADIFFAREA     0.2210 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.250 1.420 4.325 1.705 ;
        RECT  4.165 1.370 4.250 1.705 ;
        RECT  4.015 1.370 4.165 1.700 ;
        RECT  3.825 1.290 4.015 1.700 ;
        RECT  3.805 1.290 3.825 1.580 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.290 2.175 1.580 ;
        RECT  1.965 1.290 1.975 1.965 ;
        RECT  1.815 1.420 1.965 1.965 ;
        RECT  1.715 1.705 1.815 1.965 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.575 -0.250 6.900 0.250 ;
        RECT  6.315 -0.250 6.575 0.405 ;
        RECT  5.295 -0.250 6.315 0.250 ;
        RECT  5.035 -0.250 5.295 0.405 ;
        RECT  4.125 -0.250 5.035 0.250 ;
        RECT  3.865 -0.250 4.125 0.405 ;
        RECT  1.915 -0.250 3.865 0.250 ;
        RECT  1.655 -0.250 1.915 0.405 ;
        RECT  0.385 -0.250 1.655 0.250 ;
        RECT  0.125 -0.250 0.385 0.745 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 3.440 6.900 3.940 ;
        RECT  6.515 2.840 6.775 3.940 ;
        RECT  5.610 3.440 6.515 3.940 ;
        RECT  5.350 3.070 5.610 3.940 ;
        RECT  4.480 3.440 5.350 3.940 ;
        RECT  4.220 3.285 4.480 3.940 ;
        RECT  2.235 3.440 4.220 3.940 ;
        RECT  1.975 3.285 2.235 3.940 ;
        RECT  0.385 3.440 1.975 3.940 ;
        RECT  0.125 2.555 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 0.610 6.385 1.495 ;
        RECT  6.030 0.610 6.225 0.770 ;
        RECT  5.770 0.510 6.030 0.770 ;
        RECT  5.530 0.610 5.770 0.770 ;
        RECT  5.370 0.610 5.530 2.890 ;
        RECT  4.990 2.730 5.370 2.890 ;
        RECT  5.030 0.700 5.190 2.215 ;
        RECT  4.725 0.700 5.030 0.860 ;
        RECT  4.725 2.730 4.990 3.105 ;
        RECT  4.300 2.390 4.850 2.550 ;
        RECT  4.645 1.080 4.805 2.165 ;
        RECT  4.465 0.520 4.725 0.860 ;
        RECT  4.040 2.945 4.725 3.105 ;
        RECT  4.445 1.080 4.645 1.240 ;
        RECT  3.960 2.005 4.645 2.165 ;
        RECT  3.615 0.700 4.465 0.860 ;
        RECT  4.140 2.390 4.300 2.745 ;
        RECT  1.215 2.585 4.140 2.745 ;
        RECT  3.880 2.945 4.040 3.255 ;
        RECT  3.800 2.005 3.960 2.405 ;
        RECT  2.975 2.245 3.800 2.405 ;
        RECT  3.455 0.700 3.615 2.050 ;
        RECT  3.155 1.890 3.455 2.050 ;
        RECT  2.975 1.410 3.275 1.570 ;
        RECT  2.765 0.950 3.025 1.225 ;
        RECT  2.815 1.410 2.975 2.405 ;
        RECT  2.665 2.945 2.925 3.255 ;
        RECT  1.535 2.175 2.815 2.335 ;
        RECT  1.325 0.950 2.765 1.110 ;
        RECT  0.765 2.945 2.665 3.105 ;
        RECT  0.765 0.610 1.535 0.770 ;
        RECT  1.375 1.705 1.535 2.335 ;
        RECT  1.285 1.705 1.375 1.965 ;
        RECT  1.105 0.950 1.325 1.250 ;
        RECT  1.105 2.485 1.215 2.745 ;
        RECT  0.945 0.950 1.105 2.745 ;
        RECT  0.605 0.610 0.765 3.105 ;
        RECT  0.575 2.695 0.605 2.955 ;
    END
END TLATSRXL

MACRO TLATX4
    CLASS CORE ;
    FOREIGN TLATX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.025 1.700 7.235 2.400 ;
        RECT  6.795 1.700 7.025 2.395 ;
        RECT  6.775 1.055 6.795 2.395 ;
        RECT  6.725 1.055 6.775 2.585 ;
        RECT  6.555 0.695 6.725 3.010 ;
        RECT  6.465 0.695 6.555 1.295 ;
        RECT  6.465 2.070 6.555 3.010 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 1.290 5.855 2.220 ;
        RECT  5.445 0.695 5.705 2.220 ;
        END
        ANTENNADIFFAREA     0.8056 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.895 ;
        RECT  0.110 1.515 0.125 1.895 ;
        END
        ANTENNAGATEAREA     0.1573 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 1.485 1.835 1.990 ;
        RECT  1.505 1.700 1.575 1.990 ;
        END
        ANTENNAGATEAREA     0.4628 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 -0.250 7.360 0.250 ;
        RECT  6.975 -0.250 7.235 1.095 ;
        RECT  6.215 -0.250 6.975 0.250 ;
        RECT  5.955 -0.250 6.215 1.095 ;
        RECT  5.190 -0.250 5.955 0.250 ;
        RECT  4.930 -0.250 5.190 1.095 ;
        RECT  3.485 -0.250 4.930 0.250 ;
        RECT  3.225 -0.250 3.485 0.405 ;
        RECT  1.695 -0.250 3.225 0.250 ;
        RECT  1.435 -0.250 1.695 0.735 ;
        RECT  0.385 -0.250 1.435 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.235 3.440 7.360 3.940 ;
        RECT  6.975 2.600 7.235 3.940 ;
        RECT  6.215 3.440 6.975 3.940 ;
        RECT  5.955 2.940 6.215 3.940 ;
        RECT  5.165 3.440 5.955 3.940 ;
        RECT  4.905 3.285 5.165 3.940 ;
        RECT  3.415 3.440 4.905 3.940 ;
        RECT  3.155 3.285 3.415 3.940 ;
        RECT  1.580 3.440 3.155 3.940 ;
        RECT  1.320 2.955 1.580 3.940 ;
        RECT  0.385 3.440 1.320 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.260 1.580 6.360 1.840 ;
        RECT  6.100 1.580 6.260 2.760 ;
        RECT  5.225 2.600 6.100 2.760 ;
        RECT  5.065 1.275 5.225 2.760 ;
        RECT  4.750 1.275 5.065 1.440 ;
        RECT  4.705 2.600 5.065 2.760 ;
        RECT  4.405 1.620 4.885 1.780 ;
        RECT  4.610 0.655 4.750 1.440 ;
        RECT  4.545 2.250 4.705 2.940 ;
        RECT  4.590 0.550 4.610 1.440 ;
        RECT  4.350 0.550 4.590 0.815 ;
        RECT  3.270 2.780 4.545 2.940 ;
        RECT  4.365 1.110 4.405 2.050 ;
        RECT  4.245 1.110 4.365 2.600 ;
        RECT  3.985 0.655 4.350 0.815 ;
        RECT  2.585 1.110 4.245 1.270 ;
        RECT  4.205 1.890 4.245 2.600 ;
        RECT  2.560 2.440 4.205 2.600 ;
        RECT  3.940 1.480 4.065 1.640 ;
        RECT  3.725 0.470 3.985 0.815 ;
        RECT  3.780 1.480 3.940 2.260 ;
        RECT  2.315 2.100 3.780 2.260 ;
        RECT  2.795 1.760 3.585 1.920 ;
        RECT  2.635 1.465 2.795 1.920 ;
        RECT  2.535 1.465 2.635 1.745 ;
        RECT  2.375 0.685 2.585 1.285 ;
        RECT  2.435 2.440 2.560 2.775 ;
        RECT  2.175 1.465 2.535 1.625 ;
        RECT  2.400 2.440 2.435 3.215 ;
        RECT  2.175 2.615 2.400 3.215 ;
        RECT  2.325 0.685 2.375 0.945 ;
        RECT  2.215 1.805 2.315 2.260 ;
        RECT  2.055 1.805 2.215 2.335 ;
        RECT  2.015 1.140 2.175 1.625 ;
        RECT  1.605 2.175 2.055 2.335 ;
        RECT  1.265 1.140 2.015 1.300 ;
        RECT  1.445 2.175 1.605 2.775 ;
        RECT  0.785 2.615 1.445 2.775 ;
        RECT  1.255 1.140 1.265 2.400 ;
        RECT  1.105 0.525 1.255 2.400 ;
        RECT  1.095 0.525 1.105 1.300 ;
        RECT  0.925 2.140 1.105 2.400 ;
        RECT  0.925 0.525 1.095 0.785 ;
        RECT  0.710 1.640 0.925 1.900 ;
        RECT  0.710 1.035 0.815 1.295 ;
        RECT  0.710 2.615 0.785 2.910 ;
        RECT  0.550 1.035 0.710 2.910 ;
        RECT  0.525 2.650 0.550 2.910 ;
    END
END TLATX4

MACRO TLATX2
    CLASS CORE ;
    FOREIGN TLATX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.520 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.185 0.675 5.395 2.955 ;
        RECT  5.135 0.675 5.185 1.275 ;
        RECT  5.135 2.015 5.185 2.955 ;
        END
        ANTENNADIFFAREA     0.7208 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 1.290 4.475 1.765 ;
        RECT  4.275 1.290 4.375 2.895 ;
        RECT  4.115 1.210 4.275 2.895 ;
        RECT  4.100 1.210 4.115 1.370 ;
        RECT  3.840 1.010 4.100 1.370 ;
        END
        ANTENNADIFFAREA     0.7458 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 0.880 0.370 1.975 ;
        RECT  0.110 1.715 0.125 1.975 ;
        END
        ANTENNAGATEAREA     0.0858 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 1.395 1.865 1.655 ;
        RECT  1.715 1.395 1.765 1.985 ;
        RECT  1.605 1.395 1.715 1.990 ;
        RECT  1.505 1.700 1.605 1.990 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 -0.250 5.520 0.250 ;
        RECT  4.625 -0.250 4.885 0.685 ;
        RECT  3.395 -0.250 4.625 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  1.605 -0.250 3.135 0.250 ;
        RECT  1.345 -0.250 1.605 0.405 ;
        RECT  0.385 -0.250 1.345 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 3.440 5.520 3.940 ;
        RECT  4.625 2.105 4.885 3.940 ;
        RECT  3.285 3.440 4.625 3.940 ;
        RECT  3.025 3.285 3.285 3.940 ;
        RECT  1.515 3.440 3.025 3.940 ;
        RECT  1.255 2.955 1.515 3.940 ;
        RECT  0.385 3.440 1.255 3.940 ;
        RECT  0.125 2.895 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.845 1.575 5.005 1.835 ;
        RECT  4.685 0.870 4.845 1.835 ;
        RECT  4.440 0.870 4.685 1.030 ;
        RECT  4.280 0.590 4.440 1.030 ;
        RECT  3.975 0.590 4.280 0.750 ;
        RECT  3.715 0.550 3.975 0.750 ;
        RECT  3.775 1.550 3.935 2.645 ;
        RECT  3.655 1.550 3.775 1.710 ;
        RECT  3.565 2.385 3.775 2.645 ;
        RECT  3.655 0.590 3.715 0.750 ;
        RECT  3.495 0.590 3.655 1.710 ;
        RECT  2.980 1.940 3.590 2.200 ;
        RECT  3.160 1.395 3.495 1.710 ;
        RECT  2.820 0.710 2.980 2.955 ;
        RECT  2.525 0.710 2.820 0.870 ;
        RECT  2.345 2.795 2.820 2.955 ;
        RECT  2.480 1.050 2.640 2.135 ;
        RECT  2.345 2.355 2.605 2.615 ;
        RECT  2.265 0.495 2.525 0.870 ;
        RECT  1.560 1.050 2.480 1.210 ;
        RECT  2.395 1.875 2.480 2.135 ;
        RECT  2.210 2.355 2.345 2.515 ;
        RECT  2.085 2.795 2.345 3.055 ;
        RECT  2.210 1.395 2.300 1.655 ;
        RECT  2.050 1.395 2.210 2.515 ;
        RECT  1.220 2.355 2.050 2.515 ;
        RECT  1.400 0.725 1.560 1.210 ;
        RECT  0.955 0.725 1.400 0.885 ;
        RECT  1.125 1.065 1.220 2.515 ;
        RECT  1.060 1.065 1.125 2.775 ;
        RECT  0.925 1.065 1.060 1.325 ;
        RECT  0.965 2.355 1.060 2.775 ;
        RECT  0.925 2.615 0.965 2.775 ;
        RECT  0.745 0.500 0.955 0.885 ;
        RECT  0.665 2.615 0.925 3.030 ;
        RECT  0.785 1.655 0.880 1.915 ;
        RECT  0.745 1.655 0.785 2.415 ;
        RECT  0.695 0.500 0.745 2.415 ;
        RECT  0.585 0.725 0.695 2.415 ;
        RECT  0.525 2.155 0.585 2.415 ;
    END
END TLATX2

MACRO TLATX1
    CLASS CORE ;
    FOREIGN TLATX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.515 4.475 2.585 ;
        RECT  4.415 1.515 4.425 2.715 ;
        RECT  4.265 1.025 4.415 2.715 ;
        RECT  4.255 1.025 4.265 2.335 ;
        END
        ANTENNADIFFAREA     0.4247 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.915 0.680 4.075 2.680 ;
        RECT  3.595 0.680 3.915 0.840 ;
        RECT  3.805 2.335 3.915 2.680 ;
        RECT  3.565 2.520 3.805 2.680 ;
        RECT  3.335 0.580 3.595 0.840 ;
        RECT  3.345 2.520 3.565 2.855 ;
        RECT  3.305 2.595 3.345 2.855 ;
        END
        ANTENNADIFFAREA     0.3796 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.475 0.445 1.735 ;
        RECT  0.125 1.120 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0676 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.700 1.715 1.990 ;
        RECT  1.505 1.180 1.555 1.990 ;
        RECT  1.395 1.180 1.505 1.925 ;
        END
        ANTENNAGATEAREA     0.1469 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 -0.250 4.600 0.250 ;
        RECT  3.940 -0.250 4.200 0.405 ;
        RECT  3.045 -0.250 3.940 0.250 ;
        RECT  2.785 -0.250 3.045 0.405 ;
        RECT  1.465 -0.250 2.785 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 3.440 4.600 3.940 ;
        RECT  3.815 3.285 4.075 3.940 ;
        RECT  2.995 3.440 3.815 3.940 ;
        RECT  2.735 3.285 2.995 3.940 ;
        RECT  1.275 3.440 2.735 3.940 ;
        RECT  1.115 2.975 1.275 3.940 ;
        RECT  0.385 3.440 1.115 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.625 1.175 3.735 1.760 ;
        RECT  3.575 1.175 3.625 2.295 ;
        RECT  3.365 1.175 3.575 1.335 ;
        RECT  3.465 1.550 3.575 2.295 ;
        RECT  3.085 2.135 3.465 2.295 ;
        RECT  2.585 1.495 3.255 1.755 ;
        RECT  2.925 2.135 3.085 3.010 ;
        RECT  2.505 2.850 2.925 3.010 ;
        RECT  2.425 0.770 2.585 2.670 ;
        RECT  2.265 0.770 2.425 0.930 ;
        RECT  1.820 2.510 2.425 2.670 ;
        RECT  2.020 2.850 2.280 3.110 ;
        RECT  2.105 0.670 2.265 0.930 ;
        RECT  2.055 1.180 2.145 1.440 ;
        RECT  1.895 1.180 2.055 2.330 ;
        RECT  1.640 2.850 2.020 3.010 ;
        RECT  1.885 0.695 1.895 1.440 ;
        RECT  1.640 2.170 1.895 2.330 ;
        RECT  1.735 0.695 1.885 1.390 ;
        RECT  1.215 0.695 1.735 0.855 ;
        RECT  1.480 2.170 1.640 3.010 ;
        RECT  1.055 0.695 1.215 2.765 ;
        RECT  0.895 0.695 1.055 0.855 ;
        RECT  0.485 2.605 1.055 2.765 ;
        RECT  0.715 0.470 0.895 0.855 ;
        RECT  0.795 1.515 0.875 1.780 ;
        RECT  0.565 2.945 0.825 3.220 ;
        RECT  0.795 1.035 0.815 1.295 ;
        RECT  0.635 1.035 0.795 2.330 ;
        RECT  0.635 0.470 0.715 0.630 ;
        RECT  0.555 1.035 0.635 1.295 ;
        RECT  0.535 1.960 0.635 2.330 ;
        RECT  0.305 2.945 0.565 3.105 ;
        RECT  0.305 2.170 0.535 2.330 ;
        RECT  0.145 2.170 0.305 3.105 ;
    END
END TLATX1

MACRO TLATXL
    CLASS CORE ;
    FOREIGN TLATXL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.425 1.515 4.475 2.810 ;
        RECT  4.265 1.025 4.425 2.810 ;
        RECT  4.205 2.305 4.265 2.810 ;
        END
        ANTENNADIFFAREA     0.2827 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 0.595 4.085 2.100 ;
        RECT  3.925 0.595 4.020 2.855 ;
        RECT  3.680 0.595 3.925 0.755 ;
        RECT  3.860 1.940 3.925 2.855 ;
        RECT  3.805 2.110 3.860 2.855 ;
        RECT  3.190 2.595 3.805 2.855 ;
        RECT  3.420 0.495 3.680 0.755 ;
        END
        ANTENNADIFFAREA     0.2340 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.475 0.445 1.735 ;
        RECT  0.125 1.120 0.335 1.990 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 1.700 1.715 1.990 ;
        RECT  1.505 1.120 1.555 1.990 ;
        RECT  1.395 1.120 1.505 1.925 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 -0.250 4.600 0.250 ;
        RECT  4.020 -0.250 4.280 0.405 ;
        RECT  3.095 -0.250 4.020 0.250 ;
        RECT  2.835 -0.250 3.095 0.405 ;
        RECT  1.465 -0.250 2.835 0.250 ;
        RECT  1.205 -0.250 1.465 0.405 ;
        RECT  0.385 -0.250 1.205 0.250 ;
        RECT  0.125 -0.250 0.385 0.405 ;
        RECT  0.000 -0.250 0.125 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.820 3.440 4.600 3.940 ;
        RECT  3.560 3.285 3.820 3.940 ;
        RECT  2.975 3.440 3.560 3.940 ;
        RECT  2.715 3.285 2.975 3.940 ;
        RECT  1.325 3.440 2.715 3.940 ;
        RECT  1.065 2.860 1.325 3.940 ;
        RECT  0.385 3.440 1.065 3.940 ;
        RECT  0.125 3.285 0.385 3.940 ;
        RECT  0.000 3.440 0.125 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.625 1.500 3.745 1.760 ;
        RECT  3.625 1.005 3.680 1.265 ;
        RECT  3.465 1.005 3.625 2.295 ;
        RECT  3.420 1.005 3.465 1.265 ;
        RECT  3.010 2.135 3.465 2.295 ;
        RECT  2.670 1.695 3.245 1.955 ;
        RECT  2.850 2.135 3.010 3.060 ;
        RECT  2.535 2.900 2.850 3.060 ;
        RECT  2.510 0.780 2.670 2.510 ;
        RECT  2.275 2.900 2.535 3.160 ;
        RECT  2.350 0.780 2.510 0.940 ;
        RECT  2.065 2.350 2.510 2.510 ;
        RECT  2.090 0.680 2.350 0.940 ;
        RECT  2.145 1.910 2.295 2.170 ;
        RECT  1.985 1.120 2.145 2.170 ;
        RECT  1.805 2.350 2.065 2.610 ;
        RECT  1.895 1.120 1.985 1.385 ;
        RECT  1.735 0.775 1.895 1.385 ;
        RECT  1.215 0.775 1.735 0.935 ;
        RECT  1.055 0.690 1.215 2.680 ;
        RECT  0.895 0.690 1.055 0.855 ;
        RECT  0.485 2.520 1.055 2.680 ;
        RECT  0.715 0.490 0.895 0.855 ;
        RECT  0.815 1.515 0.875 1.780 ;
        RECT  0.565 2.860 0.825 3.120 ;
        RECT  0.655 1.035 0.815 2.330 ;
        RECT  0.635 0.490 0.715 0.650 ;
        RECT  0.555 1.035 0.655 1.295 ;
        RECT  0.555 1.960 0.655 2.330 ;
        RECT  0.305 2.860 0.565 3.020 ;
        RECT  0.305 2.170 0.555 2.330 ;
        RECT  0.145 2.170 0.305 3.020 ;
    END
END TLATXL

MACRO SMDFFHQX8
    CLASS CORE ;
    FOREIGN SMDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.540 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.335 6.615 1.495 ;
        RECT  5.945 0.585 6.105 1.495 ;
        RECT  3.790 0.585 5.945 0.745 ;
        RECT  3.630 0.470 3.790 0.745 ;
        RECT  1.530 0.470 3.630 0.630 ;
        RECT  1.525 0.470 1.530 0.695 ;
        RECT  1.245 0.430 1.525 0.745 ;
        RECT  1.230 0.535 1.245 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.745 7.185 1.905 ;
        RECT  5.850 1.700 5.855 1.990 ;
        RECT  5.645 1.675 5.850 1.990 ;
        RECT  5.485 1.575 5.645 1.835 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.900 1.105 21.955 2.585 ;
        RECT  21.640 0.695 21.900 2.895 ;
        RECT  21.035 1.290 21.640 1.990 ;
        RECT  20.875 1.290 21.035 2.175 ;
        RECT  20.615 0.695 20.875 2.895 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 1.185 9.640 1.680 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  10.915 1.160 11.360 1.420 ;
        RECT  10.705 1.160 10.915 1.580 ;
        RECT  10.420 1.160 10.705 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.410 -0.250 22.540 0.250 ;
        RECT  22.150 -0.250 22.410 1.115 ;
        RECT  21.385 -0.250 22.150 0.250 ;
        RECT  21.125 -0.250 21.385 1.065 ;
        RECT  20.325 -0.250 21.125 0.250 ;
        RECT  20.065 -0.250 20.325 0.405 ;
        RECT  19.445 -0.250 20.065 0.250 ;
        RECT  19.185 -0.250 19.445 0.405 ;
        RECT  16.610 -0.250 19.185 0.250 ;
        RECT  16.350 -0.250 16.610 0.785 ;
        RECT  15.530 -0.250 16.350 0.250 ;
        RECT  15.270 -0.250 15.530 0.865 ;
        RECT  14.420 -0.250 15.270 0.250 ;
        RECT  14.160 -0.250 14.420 0.405 ;
        RECT  12.690 -0.250 14.160 0.250 ;
        RECT  12.430 -0.250 12.690 0.405 ;
        RECT  11.405 -0.250 12.430 0.250 ;
        RECT  11.145 -0.250 11.405 0.405 ;
        RECT  10.325 -0.250 11.145 0.250 ;
        RECT  10.065 -0.250 10.325 0.405 ;
        RECT  9.275 -0.250 10.065 0.250 ;
        RECT  9.015 -0.250 9.275 0.405 ;
        RECT  7.375 -0.250 9.015 0.250 ;
        RECT  7.115 -0.250 7.375 0.405 ;
        RECT  6.235 -0.250 7.115 0.250 ;
        RECT  5.975 -0.250 6.235 0.405 ;
        RECT  4.235 -0.250 5.975 0.250 ;
        RECT  3.975 -0.250 4.235 0.405 ;
        RECT  0.815 -0.250 3.975 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.410 3.440 22.540 3.940 ;
        RECT  22.150 2.255 22.410 3.940 ;
        RECT  21.385 3.440 22.150 3.940 ;
        RECT  21.125 2.595 21.385 3.940 ;
        RECT  20.360 3.440 21.125 3.940 ;
        RECT  20.100 2.935 20.360 3.940 ;
        RECT  19.455 3.440 20.100 3.940 ;
        RECT  19.195 2.475 19.455 3.940 ;
        RECT  16.895 3.440 19.195 3.940 ;
        RECT  16.635 3.285 16.895 3.940 ;
        RECT  15.815 3.440 16.635 3.940 ;
        RECT  15.555 3.285 15.815 3.940 ;
        RECT  14.545 3.440 15.555 3.940 ;
        RECT  14.285 2.890 14.545 3.940 ;
        RECT  12.835 3.440 14.285 3.940 ;
        RECT  12.575 3.285 12.835 3.940 ;
        RECT  11.745 3.440 12.575 3.940 ;
        RECT  11.485 3.285 11.745 3.940 ;
        RECT  9.795 3.440 11.485 3.940 ;
        RECT  9.535 3.285 9.795 3.940 ;
        RECT  7.695 3.440 9.535 3.940 ;
        RECT  7.435 3.285 7.695 3.940 ;
        RECT  6.645 3.440 7.435 3.940 ;
        RECT  6.385 2.945 6.645 3.940 ;
        RECT  5.490 3.440 6.385 3.940 ;
        RECT  5.230 3.285 5.490 3.940 ;
        RECT  4.285 3.405 5.230 3.940 ;
        RECT  4.025 3.095 4.285 3.940 ;
        RECT  0.815 3.440 4.025 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.330 1.490 20.430 1.750 ;
        RECT  20.170 0.605 20.330 1.750 ;
        RECT  18.540 0.605 20.170 0.765 ;
        RECT  19.915 2.425 19.965 2.685 ;
        RECT  19.755 0.945 19.915 2.685 ;
        RECT  19.650 0.945 19.755 1.105 ;
        RECT  19.185 1.555 19.755 1.845 ;
        RECT  19.705 2.425 19.755 2.685 ;
        RECT  18.845 1.055 19.005 3.100 ;
        RECT  18.710 1.055 18.845 1.215 ;
        RECT  14.985 2.940 18.845 3.100 ;
        RECT  18.550 0.955 18.710 1.215 ;
        RECT  18.505 1.955 18.665 2.215 ;
        RECT  18.370 0.515 18.540 0.775 ;
        RECT  18.370 1.955 18.505 2.115 ;
        RECT  18.210 0.515 18.370 2.115 ;
        RECT  18.055 2.465 18.315 2.725 ;
        RECT  17.520 0.665 18.210 0.830 ;
        RECT  17.805 1.955 18.210 2.115 ;
        RECT  17.295 2.565 18.055 2.725 ;
        RECT  17.930 1.035 18.030 1.295 ;
        RECT  17.770 1.035 17.930 1.605 ;
        RECT  17.545 1.955 17.805 2.215 ;
        RECT  17.245 1.445 17.770 1.605 ;
        RECT  17.260 0.665 17.520 1.265 ;
        RECT  17.245 2.125 17.295 2.725 ;
        RECT  17.085 1.445 17.245 2.725 ;
        RECT  17.015 1.445 17.085 1.605 ;
        RECT  17.035 2.125 17.085 2.725 ;
        RECT  16.355 2.565 17.035 2.725 ;
        RECT  16.855 1.035 17.015 1.605 ;
        RECT  16.750 1.035 16.855 1.295 ;
        RECT  16.070 1.135 16.750 1.295 ;
        RECT  15.320 1.585 16.525 1.845 ;
        RECT  16.095 2.125 16.355 2.725 ;
        RECT  15.585 2.360 16.095 2.520 ;
        RECT  15.810 0.690 16.070 1.295 ;
        RECT  15.325 2.360 15.585 2.620 ;
        RECT  15.160 1.135 15.320 2.180 ;
        RECT  14.790 1.135 15.160 1.295 ;
        RECT  14.905 2.020 15.160 2.180 ;
        RECT  14.730 0.535 14.990 0.795 ;
        RECT  14.825 2.550 14.985 3.100 ;
        RECT  14.645 2.020 14.905 2.280 ;
        RECT  14.090 2.550 14.825 2.710 ;
        RECT  14.530 1.035 14.790 1.295 ;
        RECT  13.935 0.585 14.730 0.745 ;
        RECT  14.420 1.475 14.680 1.735 ;
        RECT  13.685 2.020 14.645 2.180 ;
        RECT  13.585 1.085 14.530 1.245 ;
        RECT  13.245 1.475 14.420 1.635 ;
        RECT  13.930 2.550 14.090 2.765 ;
        RECT  13.775 0.480 13.935 0.745 ;
        RECT  13.245 2.605 13.930 2.765 ;
        RECT  13.255 2.945 13.855 3.215 ;
        RECT  13.060 0.480 13.775 0.640 ;
        RECT  13.425 2.020 13.685 2.280 ;
        RECT  13.425 0.820 13.585 1.245 ;
        RECT  13.310 0.820 13.425 0.980 ;
        RECT  8.695 2.945 13.255 3.105 ;
        RECT  13.085 1.245 13.245 2.765 ;
        RECT  12.920 1.245 13.085 1.405 ;
        RECT  9.980 2.605 13.085 2.765 ;
        RECT  12.900 0.480 13.060 0.920 ;
        RECT  12.660 1.145 12.920 1.405 ;
        RECT  12.470 1.610 12.905 1.885 ;
        RECT  12.470 0.760 12.900 0.920 ;
        RECT  12.310 0.760 12.470 2.285 ;
        RECT  11.890 0.885 12.310 1.145 ;
        RECT  12.295 2.125 12.310 2.285 ;
        RECT  12.035 2.125 12.295 2.385 ;
        RECT  11.700 1.650 12.125 1.935 ;
        RECT  10.335 2.225 12.035 2.385 ;
        RECT  11.540 0.710 11.700 1.935 ;
        RECT  10.865 0.710 11.540 0.870 ;
        RECT  10.545 1.775 11.540 1.935 ;
        RECT  10.605 0.610 10.865 0.870 ;
        RECT  10.285 1.775 10.545 2.040 ;
        RECT  9.820 0.710 9.980 2.765 ;
        RECT  9.785 0.710 9.820 0.870 ;
        RECT  9.525 0.610 9.785 0.870 ;
        RECT  9.140 1.955 9.255 2.555 ;
        RECT  8.995 0.745 9.140 2.555 ;
        RECT  8.980 0.745 8.995 2.120 ;
        RECT  8.735 0.745 8.980 0.905 ;
        RECT  8.475 0.645 8.735 0.905 ;
        RECT  8.535 1.085 8.695 3.105 ;
        RECT  8.295 1.085 8.535 1.245 ;
        RECT  7.135 2.945 8.535 3.105 ;
        RECT  8.265 1.425 8.325 2.715 ;
        RECT  8.225 0.595 8.295 1.245 ;
        RECT  8.165 1.425 8.265 2.765 ;
        RECT  8.135 0.495 8.225 1.245 ;
        RECT  7.955 1.425 8.165 1.585 ;
        RECT  8.005 2.505 8.165 2.765 ;
        RECT  7.965 0.495 8.135 0.755 ;
        RECT  7.795 1.055 7.955 1.585 ;
        RECT  7.615 1.795 7.895 2.055 ;
        RECT  7.565 1.055 7.795 1.215 ;
        RECT  7.455 1.395 7.615 2.275 ;
        RECT  7.385 1.395 7.455 1.555 ;
        RECT  7.095 2.115 7.455 2.275 ;
        RECT  7.225 0.995 7.385 1.555 ;
        RECT  6.815 0.995 7.225 1.155 ;
        RECT  6.975 2.520 7.135 3.105 ;
        RECT  4.965 2.520 6.975 2.680 ;
        RECT  6.555 0.895 6.815 1.155 ;
        RECT  4.625 2.860 6.185 3.020 ;
        RECT  5.305 2.170 6.065 2.330 ;
        RECT  5.305 1.045 5.495 1.305 ;
        RECT  5.235 1.045 5.305 2.330 ;
        RECT  5.145 1.145 5.235 2.330 ;
        RECT  4.575 1.635 5.145 1.895 ;
        RECT  4.805 2.415 4.965 2.680 ;
        RECT  4.395 0.925 4.815 1.085 ;
        RECT  4.055 2.415 4.805 2.575 ;
        RECT  4.395 2.075 4.760 2.235 ;
        RECT  4.465 2.755 4.625 3.020 ;
        RECT  3.825 2.755 4.465 2.915 ;
        RECT  4.235 0.925 4.395 2.235 ;
        RECT  3.435 0.925 4.235 1.085 ;
        RECT  3.895 1.400 4.055 2.575 ;
        RECT  3.840 1.400 3.895 1.560 ;
        RECT  3.485 2.415 3.895 2.575 ;
        RECT  3.580 1.300 3.840 1.560 ;
        RECT  3.665 2.755 3.825 3.220 ;
        RECT  1.200 3.060 3.665 3.220 ;
        RECT  3.325 2.415 3.485 2.880 ;
        RECT  3.275 0.810 3.435 1.085 ;
        RECT  1.710 2.720 3.325 2.880 ;
        RECT  3.145 1.300 3.315 1.560 ;
        RECT  2.065 0.925 3.275 1.085 ;
        RECT  3.055 1.300 3.145 2.480 ;
        RECT  2.985 1.350 3.055 2.480 ;
        RECT  2.245 2.220 2.985 2.380 ;
        RECT  2.195 1.320 2.275 1.480 ;
        RECT  2.195 2.220 2.245 2.480 ;
        RECT  2.035 1.320 2.195 2.480 ;
        RECT  1.905 0.810 2.065 1.085 ;
        RECT  2.015 1.320 2.035 1.480 ;
        RECT  1.985 2.220 2.035 2.480 ;
        RECT  1.710 1.210 1.760 1.470 ;
        RECT  1.550 1.210 1.710 2.880 ;
        RECT  1.500 1.210 1.550 1.470 ;
        RECT  1.445 2.420 1.550 2.680 ;
        RECT  1.040 2.580 1.200 3.220 ;
        RECT  0.385 2.580 1.040 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.125 1.025 0.225 2.515 ;
        RECT  0.115 1.035 0.125 2.515 ;
    END
END SMDFFHQX8

MACRO SMDFFHQX4
    CLASS CORE ;
    FOREIGN SMDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.160 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 1.345 6.445 1.505 ;
        RECT  5.945 0.585 6.105 1.505 ;
        RECT  3.760 0.585 5.945 0.745 ;
        RECT  3.600 0.470 3.760 0.745 ;
        RECT  1.530 0.470 3.600 0.630 ;
        RECT  1.525 0.470 1.530 0.695 ;
        RECT  1.245 0.430 1.525 0.745 ;
        RECT  1.230 0.535 1.245 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.635 0.585 0.795 1.580 ;
        RECT  0.585 1.105 0.635 1.580 ;
        RECT  0.455 1.315 0.585 1.575 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 1.745 7.015 1.905 ;
        RECT  6.105 1.700 6.315 1.990 ;
        RECT  5.485 1.700 6.105 1.870 ;
        RECT  5.325 1.575 5.485 1.870 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.525 1.105 20.575 2.585 ;
        RECT  20.515 0.695 20.525 2.585 ;
        RECT  20.265 0.695 20.515 2.895 ;
        RECT  20.255 1.510 20.265 2.895 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.325 1.290 9.535 1.670 ;
        RECT  9.045 1.335 9.325 1.670 ;
        END
        ANTENNAGATEAREA     0.2730 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  10.455 1.160 10.680 1.420 ;
        RECT  10.245 1.160 10.455 1.580 ;
        RECT  10.080 1.160 10.245 1.420 ;
        END
        ANTENNAGATEAREA     0.4238 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.035 -0.250 21.160 0.250 ;
        RECT  20.775 -0.250 21.035 1.115 ;
        RECT  19.975 -0.250 20.775 0.250 ;
        RECT  19.715 -0.250 19.975 0.405 ;
        RECT  19.175 -0.250 19.715 0.250 ;
        RECT  18.915 -0.250 19.175 0.405 ;
        RECT  16.385 -0.250 18.915 0.250 ;
        RECT  16.125 -0.250 16.385 0.785 ;
        RECT  15.275 -0.250 16.125 0.250 ;
        RECT  15.015 -0.250 15.275 0.865 ;
        RECT  14.000 -0.250 15.015 0.250 ;
        RECT  13.740 -0.250 14.000 0.405 ;
        RECT  12.255 -0.250 13.740 0.250 ;
        RECT  11.995 -0.250 12.255 0.405 ;
        RECT  11.310 -0.250 11.995 0.250 ;
        RECT  11.050 -0.250 11.310 0.405 ;
        RECT  10.230 -0.250 11.050 0.250 ;
        RECT  9.970 -0.250 10.230 0.405 ;
        RECT  9.020 -0.250 9.970 0.250 ;
        RECT  8.760 -0.250 9.020 0.405 ;
        RECT  7.140 -0.250 8.760 0.250 ;
        RECT  6.880 -0.250 7.140 0.405 ;
        RECT  6.075 -0.250 6.880 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.200 -0.250 5.815 0.250 ;
        RECT  3.940 -0.250 4.200 0.405 ;
        RECT  0.815 -0.250 3.940 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.025 3.440 21.160 3.940 ;
        RECT  20.765 2.255 21.025 3.940 ;
        RECT  20.005 3.440 20.765 3.940 ;
        RECT  19.745 2.935 20.005 3.940 ;
        RECT  19.095 3.440 19.745 3.940 ;
        RECT  18.835 2.385 19.095 3.940 ;
        RECT  16.535 3.440 18.835 3.940 ;
        RECT  16.275 3.285 16.535 3.940 ;
        RECT  14.345 3.440 16.275 3.940 ;
        RECT  14.085 3.285 14.345 3.940 ;
        RECT  12.645 3.440 14.085 3.940 ;
        RECT  12.385 3.285 12.645 3.940 ;
        RECT  11.565 3.440 12.385 3.940 ;
        RECT  11.305 3.285 11.565 3.940 ;
        RECT  9.625 3.440 11.305 3.940 ;
        RECT  9.365 3.285 9.625 3.940 ;
        RECT  7.345 3.440 9.365 3.940 ;
        RECT  7.085 3.285 7.345 3.940 ;
        RECT  6.475 3.440 7.085 3.940 ;
        RECT  6.215 2.945 6.475 3.940 ;
        RECT  5.330 3.440 6.215 3.940 ;
        RECT  5.070 3.285 5.330 3.940 ;
        RECT  4.285 3.405 5.070 3.940 ;
        RECT  4.025 3.095 4.285 3.940 ;
        RECT  0.815 3.440 4.025 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.010 1.490 20.055 1.750 ;
        RECT  19.850 0.585 20.010 1.750 ;
        RECT  18.235 0.585 19.850 0.745 ;
        RECT  19.795 1.490 19.850 1.750 ;
        RECT  19.555 0.925 19.605 1.085 ;
        RECT  19.555 2.390 19.605 2.650 ;
        RECT  19.395 0.925 19.555 2.650 ;
        RECT  19.345 0.925 19.395 1.085 ;
        RECT  18.985 1.555 19.395 1.715 ;
        RECT  19.345 2.390 19.395 2.650 ;
        RECT  18.825 1.555 18.985 1.820 ;
        RECT  18.485 1.035 18.645 3.100 ;
        RECT  18.435 1.035 18.485 1.195 ;
        RECT  15.585 2.940 18.485 3.100 ;
        RECT  18.275 0.930 18.435 1.195 ;
        RECT  18.145 1.955 18.305 2.215 ;
        RECT  18.095 0.485 18.235 0.745 ;
        RECT  18.095 1.955 18.145 2.115 ;
        RECT  17.975 0.485 18.095 2.115 ;
        RECT  17.935 0.585 17.975 2.115 ;
        RECT  17.695 2.465 17.955 2.725 ;
        RECT  17.295 0.585 17.935 0.745 ;
        RECT  17.445 1.955 17.935 2.115 ;
        RECT  17.595 1.035 17.755 1.605 ;
        RECT  16.935 2.565 17.695 2.725 ;
        RECT  16.835 1.445 17.595 1.605 ;
        RECT  17.185 1.955 17.445 2.215 ;
        RECT  17.035 0.585 17.295 1.265 ;
        RECT  16.835 2.125 16.935 2.725 ;
        RECT  16.675 1.035 16.835 2.725 ;
        RECT  15.845 1.035 16.675 1.295 ;
        RECT  15.995 2.565 16.675 2.725 ;
        RECT  14.940 1.585 16.120 1.845 ;
        RECT  15.735 2.125 15.995 2.725 ;
        RECT  15.585 0.690 15.845 1.295 ;
        RECT  15.155 2.565 15.735 2.725 ;
        RECT  15.425 2.940 15.585 3.190 ;
        RECT  14.715 3.030 15.425 3.190 ;
        RECT  14.945 2.565 15.155 2.850 ;
        RECT  14.895 2.690 14.945 2.850 ;
        RECT  14.780 1.135 14.940 2.180 ;
        RECT  14.565 1.135 14.780 1.295 ;
        RECT  14.665 2.020 14.780 2.180 ;
        RECT  14.505 0.535 14.765 0.795 ;
        RECT  14.665 2.605 14.715 2.765 ;
        RECT  14.555 2.945 14.715 3.190 ;
        RECT  14.505 2.020 14.665 2.765 ;
        RECT  14.305 1.035 14.565 1.295 ;
        RECT  14.005 2.945 14.555 3.105 ;
        RECT  13.475 0.585 14.505 0.745 ;
        RECT  13.495 2.020 14.505 2.180 ;
        RECT  14.455 2.605 14.505 2.765 ;
        RECT  14.195 1.475 14.455 1.735 ;
        RECT  14.265 1.035 14.305 1.195 ;
        RECT  14.105 0.925 14.265 1.195 ;
        RECT  13.045 1.475 14.195 1.635 ;
        RECT  13.135 0.925 14.105 1.085 ;
        RECT  13.845 2.605 14.005 3.105 ;
        RECT  13.045 2.605 13.845 2.765 ;
        RECT  13.065 2.945 13.665 3.215 ;
        RECT  13.235 2.020 13.495 2.280 ;
        RECT  13.315 0.485 13.475 0.745 ;
        RECT  12.595 0.485 13.315 0.645 ;
        RECT  12.875 0.825 13.135 1.085 ;
        RECT  8.525 2.945 13.065 3.105 ;
        RECT  12.885 1.285 13.045 2.765 ;
        RECT  12.435 1.285 12.885 1.445 ;
        RECT  9.875 2.605 12.885 2.765 ;
        RECT  12.105 1.625 12.705 1.885 ;
        RECT  12.435 0.485 12.595 0.745 ;
        RECT  12.095 0.585 12.435 0.745 ;
        RECT  12.275 1.145 12.435 1.445 ;
        RECT  12.095 1.625 12.105 2.385 ;
        RECT  11.935 0.585 12.095 2.385 ;
        RECT  11.455 0.885 11.935 1.145 ;
        RECT  11.845 2.125 11.935 2.385 ;
        RECT  10.165 2.225 11.845 2.385 ;
        RECT  11.080 1.650 11.755 1.935 ;
        RECT  10.920 0.710 11.080 1.935 ;
        RECT  10.770 0.710 10.920 0.870 ;
        RECT  10.215 1.775 10.920 1.935 ;
        RECT  10.510 0.610 10.770 0.870 ;
        RECT  10.055 1.775 10.215 2.040 ;
        RECT  9.715 0.710 9.875 2.765 ;
        RECT  9.690 0.710 9.715 0.870 ;
        RECT  9.430 0.610 9.690 0.870 ;
        RECT  8.865 1.955 9.085 2.555 ;
        RECT  8.825 0.675 8.865 2.555 ;
        RECT  8.705 0.675 8.825 2.120 ;
        RECT  8.480 0.675 8.705 0.835 ;
        RECT  8.365 1.015 8.525 3.105 ;
        RECT  8.220 0.575 8.480 0.835 ;
        RECT  8.040 1.015 8.365 1.175 ;
        RECT  6.830 2.945 8.365 3.105 ;
        RECT  7.970 0.595 8.040 1.175 ;
        RECT  7.880 0.495 7.970 1.175 ;
        RECT  7.765 1.360 7.925 2.765 ;
        RECT  7.710 0.495 7.880 0.755 ;
        RECT  7.695 1.360 7.765 1.520 ;
        RECT  7.665 2.505 7.765 2.765 ;
        RECT  7.535 1.055 7.695 1.520 ;
        RECT  7.310 1.055 7.535 1.215 ;
        RECT  7.355 1.695 7.445 2.055 ;
        RECT  7.195 1.400 7.355 2.275 ;
        RECT  6.800 1.400 7.195 1.560 ;
        RECT  6.925 2.115 7.195 2.275 ;
        RECT  6.670 2.520 6.830 3.105 ;
        RECT  6.640 0.995 6.800 1.560 ;
        RECT  4.965 2.520 6.670 2.680 ;
        RECT  6.535 0.995 6.640 1.155 ;
        RECT  6.535 0.490 6.585 0.750 ;
        RECT  6.375 0.490 6.535 1.155 ;
        RECT  6.325 0.490 6.375 0.750 ;
        RECT  4.625 2.860 6.030 3.020 ;
        RECT  5.800 2.170 5.905 2.330 ;
        RECT  5.640 2.055 5.800 2.330 ;
        RECT  5.140 2.055 5.640 2.215 ;
        RECT  5.140 1.045 5.335 1.305 ;
        RECT  5.075 1.045 5.140 2.215 ;
        RECT  4.980 1.145 5.075 2.215 ;
        RECT  4.415 1.635 4.980 1.895 ;
        RECT  4.805 2.415 4.965 2.680 ;
        RECT  3.740 2.415 4.805 2.575 ;
        RECT  4.225 0.925 4.780 1.085 ;
        RECT  4.225 2.075 4.760 2.235 ;
        RECT  4.465 2.755 4.625 3.020 ;
        RECT  3.825 2.755 4.465 2.915 ;
        RECT  4.065 0.925 4.225 2.235 ;
        RECT  3.420 0.925 4.065 1.085 ;
        RECT  3.740 1.300 3.840 1.560 ;
        RECT  3.665 2.755 3.825 3.220 ;
        RECT  3.580 1.300 3.740 2.575 ;
        RECT  1.200 3.060 3.665 3.220 ;
        RECT  3.485 2.415 3.580 2.575 ;
        RECT  3.325 2.415 3.485 2.880 ;
        RECT  3.260 0.810 3.420 1.085 ;
        RECT  1.710 2.720 3.325 2.880 ;
        RECT  3.145 1.300 3.315 1.560 ;
        RECT  2.065 0.925 3.260 1.085 ;
        RECT  3.055 1.300 3.145 2.480 ;
        RECT  2.985 1.350 3.055 2.480 ;
        RECT  2.245 2.220 2.985 2.380 ;
        RECT  2.175 1.320 2.275 1.480 ;
        RECT  2.175 2.220 2.245 2.480 ;
        RECT  2.015 1.320 2.175 2.480 ;
        RECT  1.905 0.810 2.065 1.085 ;
        RECT  1.985 2.220 2.015 2.480 ;
        RECT  1.710 1.210 1.760 1.470 ;
        RECT  1.550 1.210 1.710 2.880 ;
        RECT  1.500 1.210 1.550 1.470 ;
        RECT  1.445 2.420 1.550 2.680 ;
        RECT  1.040 2.580 1.200 3.220 ;
        RECT  0.385 2.580 1.040 2.740 ;
        RECT  0.275 0.875 0.385 1.135 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 0.875 0.275 2.740 ;
        RECT  0.115 0.875 0.225 2.515 ;
    END
END SMDFFHQX4

MACRO SMDFFHQX2
    CLASS CORE ;
    FOREIGN SMDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.640 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.115 1.335 5.450 1.495 ;
        RECT  4.955 0.935 5.115 1.495 ;
        RECT  4.520 0.935 4.955 1.095 ;
        RECT  4.360 0.620 4.520 1.095 ;
        RECT  2.955 0.620 4.360 0.780 ;
        RECT  2.795 0.490 2.955 0.780 ;
        RECT  2.500 0.490 2.795 0.650 ;
        RECT  2.340 0.430 2.500 0.650 ;
        RECT  1.675 0.430 2.340 0.590 ;
        RECT  1.515 0.430 1.675 0.785 ;
        RECT  0.795 0.625 1.515 0.785 ;
        RECT  0.715 0.625 0.795 1.680 ;
        RECT  0.635 0.625 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.935 1.725 5.930 1.885 ;
        RECT  4.930 1.700 4.935 1.990 ;
        RECT  4.725 1.675 4.930 1.990 ;
        RECT  4.285 1.675 4.725 1.835 ;
        RECT  4.125 1.575 4.285 1.835 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.255 0.695 15.515 2.895 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.260 1.290 8.615 1.580 ;
        RECT  8.000 1.290 8.260 1.610 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.530 1.290 9.535 1.580 ;
        RECT  9.135 1.290 9.530 1.600 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 -0.250 15.640 0.250 ;
        RECT  14.715 -0.250 14.975 0.405 ;
        RECT  14.175 -0.250 14.715 0.250 ;
        RECT  13.915 -0.250 14.175 0.405 ;
        RECT  12.055 -0.250 13.915 0.250 ;
        RECT  11.795 -0.250 12.055 0.755 ;
        RECT  10.405 -0.250 11.795 0.250 ;
        RECT  10.145 -0.250 10.405 0.405 ;
        RECT  8.800 -0.250 10.145 0.250 ;
        RECT  7.780 -0.250 8.800 0.405 ;
        RECT  6.140 -0.250 7.780 0.250 ;
        RECT  5.880 -0.250 6.140 0.405 ;
        RECT  4.990 -0.250 5.880 0.250 ;
        RECT  4.730 -0.250 4.990 0.745 ;
        RECT  3.395 -0.250 4.730 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 3.440 15.640 3.940 ;
        RECT  14.715 2.890 14.975 3.940 ;
        RECT  14.125 3.440 14.715 3.940 ;
        RECT  13.865 2.890 14.125 3.940 ;
        RECT  12.195 3.440 13.865 3.940 ;
        RECT  11.935 3.285 12.195 3.940 ;
        RECT  10.435 3.440 11.935 3.940 ;
        RECT  10.175 3.285 10.435 3.940 ;
        RECT  8.415 3.440 10.175 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  6.485 3.440 8.155 3.940 ;
        RECT  6.225 3.285 6.485 3.940 ;
        RECT  5.250 3.440 6.225 3.940 ;
        RECT  4.990 2.925 5.250 3.940 ;
        RECT  4.165 3.440 4.990 3.940 ;
        RECT  3.905 3.285 4.165 3.940 ;
        RECT  3.235 3.440 3.905 3.940 ;
        RECT  3.075 3.035 3.235 3.940 ;
        RECT  0.815 3.440 3.075 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.555 2.105 14.605 2.365 ;
        RECT  14.395 1.035 14.555 2.365 ;
        RECT  14.345 2.005 14.395 2.365 ;
        RECT  13.875 2.005 14.345 2.165 ;
        RECT  14.055 0.585 14.215 1.665 ;
        RECT  13.105 0.585 14.055 0.745 ;
        RECT  13.715 1.885 13.875 2.165 ;
        RECT  13.535 2.920 13.615 3.180 ;
        RECT  13.375 0.925 13.535 3.180 ;
        RECT  13.265 0.925 13.375 1.190 ;
        RECT  13.355 2.860 13.375 3.180 ;
        RECT  11.510 2.860 13.355 3.020 ;
        RECT  13.085 1.440 13.195 2.555 ;
        RECT  13.085 0.535 13.105 0.795 ;
        RECT  13.035 0.535 13.085 2.555 ;
        RECT  12.925 0.535 13.035 1.600 ;
        RECT  12.845 0.535 12.925 0.795 ;
        RECT  12.595 1.085 12.735 2.675 ;
        RECT  12.575 0.985 12.595 2.675 ;
        RECT  12.335 0.985 12.575 1.245 ;
        RECT  12.475 2.075 12.575 2.675 ;
        RECT  11.965 2.515 12.475 2.675 ;
        RECT  12.120 1.585 12.345 1.845 ;
        RECT  11.960 1.025 12.120 2.230 ;
        RECT  11.705 2.415 11.965 2.675 ;
        RECT  11.315 1.025 11.960 1.185 ;
        RECT  11.025 2.070 11.960 2.230 ;
        RECT  10.215 0.585 11.515 0.745 ;
        RECT  11.350 2.605 11.510 3.020 ;
        RECT  10.845 1.615 11.485 1.875 ;
        RECT  10.845 2.605 11.350 2.765 ;
        RECT  11.055 0.925 11.315 1.185 ;
        RECT  11.020 3.100 11.115 3.260 ;
        RECT  10.855 2.945 11.020 3.260 ;
        RECT  7.435 2.945 10.855 3.105 ;
        RECT  10.685 1.270 10.845 2.765 ;
        RECT  10.555 1.270 10.685 1.430 ;
        RECT  8.775 2.605 10.685 2.765 ;
        RECT  10.395 1.170 10.555 1.430 ;
        RECT  10.215 1.650 10.505 1.910 ;
        RECT  10.055 0.585 10.215 2.385 ;
        RECT  9.865 0.585 10.055 0.770 ;
        RECT  8.955 2.225 10.055 2.385 ;
        RECT  9.715 0.950 9.875 1.940 ;
        RECT  9.605 0.510 9.865 0.770 ;
        RECT  9.300 0.950 9.715 1.110 ;
        RECT  9.295 1.780 9.715 1.940 ;
        RECT  9.140 0.840 9.300 1.110 ;
        RECT  9.135 1.780 9.295 2.040 ;
        RECT  8.795 0.940 8.955 1.920 ;
        RECT  8.400 0.940 8.795 1.100 ;
        RECT  8.775 1.760 8.795 1.920 ;
        RECT  8.615 1.760 8.775 2.765 ;
        RECT  8.140 0.840 8.400 1.100 ;
        RECT  7.775 1.955 7.995 2.555 ;
        RECT  7.735 0.670 7.775 2.555 ;
        RECT  7.615 0.670 7.735 2.120 ;
        RECT  7.230 0.670 7.615 0.830 ;
        RECT  7.275 1.085 7.435 3.105 ;
        RECT  7.050 1.085 7.275 1.245 ;
        RECT  6.095 2.945 7.275 3.105 ;
        RECT  6.905 1.425 7.065 2.765 ;
        RECT  6.890 0.455 7.050 1.245 ;
        RECT  6.710 1.425 6.905 1.585 ;
        RECT  6.745 2.505 6.905 2.765 ;
        RECT  6.690 0.455 6.890 0.715 ;
        RECT  6.550 1.015 6.710 1.585 ;
        RECT  6.270 1.795 6.635 2.055 ;
        RECT  6.310 1.015 6.550 1.175 ;
        RECT  6.130 1.380 6.270 2.225 ;
        RECT  6.110 0.995 6.130 2.225 ;
        RECT  5.970 0.995 6.110 1.540 ;
        RECT  6.100 2.065 6.110 2.225 ;
        RECT  5.840 2.065 6.100 2.325 ;
        RECT  5.935 2.520 6.095 3.105 ;
        RECT  5.560 0.995 5.970 1.155 ;
        RECT  3.915 2.520 5.935 2.680 ;
        RECT  5.300 0.895 5.560 1.155 ;
        RECT  4.550 2.860 4.810 3.120 ;
        RECT  4.255 2.170 4.680 2.330 ;
        RECT  3.575 2.860 4.550 3.020 ;
        RECT  4.095 2.015 4.255 2.330 ;
        RECT  3.940 1.045 4.110 1.305 ;
        RECT  3.940 2.015 4.095 2.175 ;
        RECT  3.780 1.045 3.940 2.175 ;
        RECT  3.755 2.355 3.915 2.680 ;
        RECT  3.585 1.575 3.780 1.835 ;
        RECT  2.555 2.355 3.755 2.515 ;
        RECT  3.340 1.045 3.600 1.305 ;
        RECT  3.120 2.015 3.595 2.175 ;
        RECT  3.415 2.695 3.575 3.020 ;
        RECT  2.895 2.695 3.415 2.855 ;
        RECT  3.120 1.095 3.340 1.305 ;
        RECT  2.960 1.095 3.120 2.175 ;
        RECT  2.615 1.095 2.960 1.255 ;
        RECT  2.735 2.695 2.895 3.135 ;
        RECT  1.365 2.975 2.735 3.135 ;
        RECT  2.455 0.835 2.615 1.255 ;
        RECT  2.395 2.355 2.555 2.735 ;
        RECT  2.115 0.835 2.455 0.995 ;
        RECT  1.705 2.575 2.395 2.735 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.130 2.215 2.390 ;
        RECT  1.855 0.770 2.115 0.995 ;
        RECT  1.955 1.175 2.115 2.390 ;
        RECT  1.705 1.210 1.725 1.470 ;
        RECT  1.545 1.210 1.705 2.735 ;
        RECT  1.515 1.210 1.545 2.390 ;
        RECT  1.465 1.210 1.515 1.470 ;
        RECT  1.445 2.130 1.515 2.390 ;
        RECT  1.205 2.580 1.365 3.135 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.515 ;
    END
END SMDFFHQX2

MACRO SMDFFHQX1
    CLASS CORE ;
    FOREIGN SMDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.260 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 1.385 4.900 1.545 ;
        RECT  4.200 0.585 4.360 1.545 ;
        RECT  2.955 0.585 4.200 0.745 ;
        RECT  2.795 0.470 2.955 0.745 ;
        RECT  2.460 0.470 2.795 0.630 ;
        RECT  2.300 0.465 2.460 0.630 ;
        RECT  1.645 0.465 2.300 0.625 ;
        RECT  1.485 0.465 1.645 0.805 ;
        RECT  1.305 0.645 1.485 0.805 ;
        RECT  1.145 0.645 1.305 1.380 ;
        RECT  1.045 1.105 1.145 1.380 ;
        RECT  0.795 1.220 1.045 1.380 ;
        RECT  0.770 1.220 0.795 1.580 ;
        RECT  0.715 1.220 0.770 1.680 ;
        RECT  0.610 1.220 0.715 1.730 ;
        RECT  0.585 1.290 0.610 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1170 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.725 5.380 1.885 ;
        RECT  3.975 1.700 4.015 1.990 ;
        RECT  3.815 1.660 3.975 1.990 ;
        RECT  3.805 1.700 3.815 1.990 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.025 1.105 14.135 2.175 ;
        RECT  13.865 0.695 14.025 2.680 ;
        RECT  13.565 0.695 13.865 0.855 ;
        RECT  13.675 2.520 13.865 2.680 ;
        RECT  13.505 2.520 13.675 2.995 ;
        RECT  13.305 0.595 13.565 0.855 ;
        RECT  13.245 2.520 13.505 3.165 ;
        END
        ANTENNADIFFAREA     0.3808 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.0923 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 0.880 7.235 1.620 ;
        RECT  7.025 0.880 7.040 1.170 ;
        END
        ANTENNAGATEAREA     0.0884 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.755 1.290 8.155 1.620 ;
        END
        ANTENNAGATEAREA     0.1261 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.025 -0.250 14.260 0.250 ;
        RECT  12.765 -0.250 13.025 0.405 ;
        RECT  10.970 -0.250 12.765 0.250 ;
        RECT  10.710 -0.250 10.970 0.405 ;
        RECT  9.290 -0.250 10.710 0.250 ;
        RECT  9.030 -0.250 9.290 0.405 ;
        RECT  7.340 -0.250 9.030 0.250 ;
        RECT  7.080 -0.250 7.340 0.405 ;
        RECT  5.530 -0.250 7.080 0.250 ;
        RECT  5.270 -0.250 5.530 0.405 ;
        RECT  4.515 -0.250 5.270 0.250 ;
        RECT  4.255 -0.250 4.515 0.405 ;
        RECT  3.395 -0.250 4.255 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.985 3.440 14.260 3.940 ;
        RECT  12.725 2.615 12.985 3.940 ;
        RECT  11.160 3.440 12.725 3.940 ;
        RECT  10.900 3.285 11.160 3.940 ;
        RECT  9.400 3.440 10.900 3.940 ;
        RECT  9.140 3.285 9.400 3.940 ;
        RECT  7.480 3.440 9.140 3.940 ;
        RECT  7.220 3.285 7.480 3.940 ;
        RECT  5.540 3.440 7.220 3.940 ;
        RECT  5.280 3.285 5.540 3.940 ;
        RECT  4.775 3.440 5.280 3.940 ;
        RECT  4.515 2.925 4.775 3.940 ;
        RECT  3.765 3.440 4.515 3.940 ;
        RECT  3.505 3.285 3.765 3.940 ;
        RECT  2.615 3.440 3.505 3.940 ;
        RECT  2.355 3.115 2.615 3.940 ;
        RECT  0.815 3.440 2.355 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.535 1.105 13.645 2.165 ;
        RECT  13.485 1.105 13.535 2.285 ;
        RECT  13.385 1.105 13.485 1.365 ;
        RECT  13.275 2.005 13.485 2.285 ;
        RECT  13.205 1.560 13.305 1.820 ;
        RECT  12.725 2.005 13.275 2.165 ;
        RECT  13.045 1.310 13.205 1.820 ;
        RECT  12.725 1.310 13.045 1.470 ;
        RECT  12.565 0.745 12.725 1.470 ;
        RECT  12.565 1.785 12.725 2.165 ;
        RECT  12.045 0.745 12.565 0.905 ;
        RECT  12.225 1.085 12.385 3.215 ;
        RECT  11.595 3.055 12.225 3.215 ;
        RECT  11.885 0.745 12.045 2.795 ;
        RECT  11.770 0.975 11.885 1.235 ;
        RECT  11.640 0.570 11.690 0.730 ;
        RECT  11.430 0.570 11.640 0.745 ;
        RECT  11.435 2.940 11.595 3.215 ;
        RECT  11.560 2.135 11.585 2.760 ;
        RECT  11.400 1.035 11.560 2.760 ;
        RECT  10.280 2.940 11.435 3.100 ;
        RECT  8.850 0.585 11.430 0.745 ;
        RECT  11.260 1.035 11.400 1.295 ;
        RECT  11.325 2.135 11.400 2.760 ;
        RECT  10.530 2.600 11.325 2.760 ;
        RECT  10.785 1.635 11.220 1.895 ;
        RECT  10.625 1.025 10.785 2.420 ;
        RECT  10.180 1.025 10.625 1.185 ;
        RECT  9.850 2.260 10.625 2.420 ;
        RECT  9.845 1.635 10.310 1.895 ;
        RECT  10.120 2.605 10.280 3.100 ;
        RECT  10.020 0.925 10.180 1.185 ;
        RECT  9.670 2.605 10.120 2.765 ;
        RECT  8.755 2.945 9.940 3.105 ;
        RECT  9.840 1.635 9.845 2.065 ;
        RECT  9.680 1.135 9.840 2.065 ;
        RECT  9.450 1.135 9.680 1.295 ;
        RECT  9.670 1.905 9.680 2.065 ;
        RECT  9.510 1.905 9.670 2.765 ;
        RECT  8.340 2.605 9.510 2.765 ;
        RECT  8.850 1.565 9.500 1.725 ;
        RECT  9.290 1.035 9.450 1.295 ;
        RECT  8.710 0.585 8.850 2.405 ;
        RECT  8.595 2.945 8.755 3.135 ;
        RECT  8.690 0.510 8.710 2.405 ;
        RECT  8.450 0.510 8.690 0.770 ;
        RECT  7.910 2.245 8.690 2.405 ;
        RECT  7.820 2.975 8.595 3.135 ;
        RECT  8.335 0.950 8.495 2.035 ;
        RECT  8.080 2.605 8.340 2.775 ;
        RECT  8.270 0.950 8.335 1.110 ;
        RECT  7.800 1.875 8.335 2.035 ;
        RECT  8.110 0.440 8.270 1.110 ;
        RECT  7.670 0.440 8.110 0.600 ;
        RECT  7.575 2.605 8.080 2.765 ;
        RECT  7.575 0.950 7.930 1.110 ;
        RECT  7.660 2.945 7.820 3.135 ;
        RECT  6.520 2.945 7.660 3.105 ;
        RECT  7.415 0.950 7.575 2.765 ;
        RECT  6.860 2.170 7.080 2.430 ;
        RECT  6.845 1.350 6.860 2.430 ;
        RECT  6.820 0.905 6.845 2.430 ;
        RECT  6.700 0.905 6.820 2.380 ;
        RECT  6.685 0.905 6.700 1.510 ;
        RECT  6.505 2.140 6.520 3.105 ;
        RECT  6.345 0.545 6.505 3.105 ;
        RECT  6.325 0.545 6.345 0.705 ;
        RECT  5.115 2.945 6.345 3.105 ;
        RECT  6.065 0.445 6.325 0.705 ;
        RECT  6.060 1.015 6.150 2.715 ;
        RECT  5.990 1.015 6.060 2.765 ;
        RECT  5.850 1.015 5.990 1.175 ;
        RECT  5.960 1.850 5.990 2.110 ;
        RECT  5.800 2.505 5.990 2.765 ;
        RECT  5.720 1.370 5.810 1.630 ;
        RECT  5.670 1.370 5.720 2.225 ;
        RECT  5.560 1.045 5.670 2.225 ;
        RECT  5.510 1.045 5.560 1.540 ;
        RECT  5.485 2.065 5.560 2.225 ;
        RECT  5.100 1.045 5.510 1.205 ;
        RECT  5.225 2.065 5.485 2.325 ;
        RECT  4.955 2.510 5.115 3.105 ;
        RECT  4.840 0.945 5.100 1.205 ;
        RECT  3.295 2.510 4.955 2.670 ;
        RECT  4.075 2.850 4.335 3.110 ;
        RECT  3.625 2.170 4.195 2.330 ;
        RECT  2.955 2.850 4.075 3.010 ;
        RECT  3.625 0.965 3.765 1.225 ;
        RECT  3.465 0.965 3.625 2.330 ;
        RECT  3.155 1.635 3.465 1.895 ;
        RECT  3.135 2.435 3.295 2.670 ;
        RECT  2.975 1.125 3.255 1.385 ;
        RECT  2.975 2.095 3.255 2.255 ;
        RECT  1.705 2.435 3.135 2.595 ;
        RECT  2.815 1.125 2.975 2.255 ;
        RECT  2.795 2.775 2.955 3.010 ;
        RECT  2.615 1.125 2.815 1.285 ;
        RECT  1.365 2.775 2.795 2.935 ;
        RECT  2.455 0.810 2.615 1.285 ;
        RECT  2.105 0.810 2.455 0.970 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.095 2.215 2.255 ;
        RECT  1.955 1.175 2.115 2.255 ;
        RECT  1.845 0.805 2.105 0.970 ;
        RECT  1.675 2.150 1.705 2.595 ;
        RECT  1.545 1.035 1.675 2.595 ;
        RECT  1.515 1.035 1.545 2.410 ;
        RECT  1.445 2.150 1.515 2.410 ;
        RECT  1.205 2.580 1.365 2.935 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.125 1.025 0.225 2.520 ;
        RECT  0.115 1.035 0.125 2.520 ;
    END
END SMDFFHQX1

MACRO SEDFFHQX8
    CLASS CORE ;
    FOREIGN SEDFFHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.620 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.990 1.255 2.400 ;
        RECT  0.975 1.565 1.235 2.400 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.335 6.305 1.495 ;
        RECT  5.740 1.105 5.855 1.495 ;
        RECT  5.580 0.650 5.740 1.495 ;
        RECT  4.415 0.650 5.580 0.810 ;
        RECT  4.255 0.470 4.415 0.810 ;
        RECT  1.505 0.470 4.255 0.630 ;
        RECT  1.435 0.430 1.505 0.630 ;
        RECT  1.230 0.430 1.435 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.955 1.515 21.035 1.765 ;
        RECT  20.695 0.695 20.955 2.895 ;
        RECT  19.930 1.290 20.695 1.990 ;
        RECT  19.670 0.695 19.930 2.920 ;
        END
        ANTENNADIFFAREA     1.5960 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.725 6.770 1.885 ;
        RECT  5.645 1.700 5.855 1.990 ;
        RECT  5.335 1.700 5.645 1.860 ;
        RECT  5.175 1.575 5.335 1.860 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 1.290 9.995 1.580 ;
        RECT  9.815 1.155 9.975 1.580 ;
        RECT  9.585 1.290 9.815 1.580 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.465 -0.250 21.620 0.250 ;
        RECT  21.205 -0.250 21.465 1.115 ;
        RECT  20.440 -0.250 21.205 0.250 ;
        RECT  20.180 -0.250 20.440 0.940 ;
        RECT  19.415 -0.250 20.180 0.250 ;
        RECT  19.155 -0.250 19.415 1.295 ;
        RECT  18.630 -0.250 19.155 0.250 ;
        RECT  18.370 -0.250 18.630 0.405 ;
        RECT  9.835 -0.250 18.370 0.250 ;
        RECT  9.575 -0.250 9.835 0.405 ;
        RECT  8.785 -0.250 9.575 0.250 ;
        RECT  8.525 -0.250 8.785 0.405 ;
        RECT  7.095 -0.250 8.525 0.250 ;
        RECT  6.835 -0.250 7.095 0.405 ;
        RECT  6.075 -0.250 6.835 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.855 -0.250 5.815 0.250 ;
        RECT  4.595 -0.250 4.855 0.405 ;
        RECT  0.815 -0.250 4.595 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.465 3.440 21.620 3.940 ;
        RECT  21.205 2.255 21.465 3.940 ;
        RECT  20.440 3.440 21.205 3.940 ;
        RECT  20.180 2.255 20.440 3.940 ;
        RECT  19.385 3.440 20.180 3.940 ;
        RECT  19.125 3.285 19.385 3.940 ;
        RECT  18.505 3.440 19.125 3.940 ;
        RECT  18.245 3.285 18.505 3.940 ;
        RECT  15.910 3.440 18.245 3.940 ;
        RECT  15.650 3.285 15.910 3.940 ;
        RECT  14.795 3.440 15.650 3.940 ;
        RECT  14.535 3.285 14.795 3.940 ;
        RECT  13.520 3.440 14.535 3.940 ;
        RECT  13.260 3.285 13.520 3.940 ;
        RECT  11.790 3.440 13.260 3.940 ;
        RECT  11.530 3.285 11.790 3.940 ;
        RECT  10.710 3.440 11.530 3.940 ;
        RECT  10.450 3.285 10.710 3.940 ;
        RECT  8.725 3.440 10.450 3.940 ;
        RECT  8.465 3.285 8.725 3.940 ;
        RECT  6.965 3.440 8.465 3.940 ;
        RECT  6.705 3.285 6.965 3.940 ;
        RECT  6.110 3.440 6.705 3.940 ;
        RECT  5.850 2.945 6.110 3.940 ;
        RECT  5.100 3.440 5.850 3.940 ;
        RECT  4.840 3.285 5.100 3.940 ;
        RECT  4.360 3.405 4.840 3.940 ;
        RECT  4.100 3.095 4.360 3.940 ;
        RECT  0.870 3.440 4.100 3.940 ;
        RECT  0.610 2.925 0.870 3.940 ;
        RECT  0.000 3.440 0.610 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.895 2.575 18.935 2.835 ;
        RECT  18.735 0.845 18.895 2.835 ;
        RECT  18.625 0.845 18.735 1.225 ;
        RECT  18.640 1.885 18.735 2.145 ;
        RECT  18.675 2.575 18.735 2.835 ;
        RECT  18.190 0.845 18.625 1.005 ;
        RECT  18.445 1.405 18.555 1.665 ;
        RECT  18.285 1.185 18.445 2.880 ;
        RECT  17.850 1.185 18.285 1.345 ;
        RECT  16.820 2.720 18.285 2.880 ;
        RECT  18.030 0.470 18.190 1.005 ;
        RECT  17.945 1.530 18.105 2.535 ;
        RECT  14.490 0.470 18.030 0.630 ;
        RECT  17.510 1.530 17.945 1.690 ;
        RECT  17.360 2.375 17.945 2.535 ;
        RECT  17.690 0.910 17.850 1.345 ;
        RECT  17.605 1.875 17.765 2.190 ;
        RECT  17.360 0.910 17.690 1.070 ;
        RECT  17.170 1.875 17.605 2.035 ;
        RECT  17.335 3.060 17.595 3.260 ;
        RECT  17.350 1.250 17.510 1.690 ;
        RECT  17.100 0.810 17.360 1.070 ;
        RECT  17.200 2.220 17.360 2.535 ;
        RECT  16.820 1.250 17.350 1.410 ;
        RECT  16.250 3.060 17.335 3.220 ;
        RECT  16.820 2.220 17.200 2.380 ;
        RECT  17.010 1.635 17.170 2.035 ;
        RECT  16.230 0.810 17.100 0.970 ;
        RECT  15.540 1.635 17.010 1.795 ;
        RECT  16.560 1.155 16.820 1.410 ;
        RECT  16.560 2.120 16.820 2.380 ;
        RECT  16.660 2.565 16.820 2.880 ;
        RECT  16.280 2.565 16.660 2.725 ;
        RECT  15.880 1.250 16.560 1.410 ;
        RECT  15.370 2.120 16.560 2.280 ;
        RECT  16.020 2.465 16.280 2.725 ;
        RECT  16.090 2.940 16.250 3.220 ;
        RECT  16.070 0.810 16.230 1.070 ;
        RECT  14.160 2.940 16.090 3.100 ;
        RECT  15.720 0.910 15.880 1.410 ;
        RECT  15.370 0.910 15.720 1.070 ;
        RECT  15.380 1.250 15.540 1.795 ;
        RECT  14.760 1.250 15.380 1.410 ;
        RECT  15.110 0.810 15.370 1.070 ;
        RECT  15.110 2.120 15.370 2.760 ;
        RECT  14.940 1.635 15.200 1.850 ;
        RECT  14.340 2.600 15.110 2.760 ;
        RECT  13.955 1.690 14.940 1.850 ;
        RECT  14.600 0.810 14.760 1.410 ;
        RECT  14.145 0.810 14.600 0.970 ;
        RECT  14.330 0.430 14.490 0.630 ;
        RECT  13.695 0.430 14.330 0.590 ;
        RECT  14.000 2.605 14.160 3.100 ;
        RECT  13.885 0.770 14.145 0.970 ;
        RECT  12.195 2.605 14.000 2.765 ;
        RECT  13.875 1.150 13.955 2.320 ;
        RECT  11.425 0.810 13.885 0.970 ;
        RECT  13.795 1.150 13.875 2.425 ;
        RECT  12.435 1.150 13.795 1.310 ;
        RECT  13.615 2.160 13.795 2.425 ;
        RECT  13.535 0.430 13.695 0.630 ;
        RECT  12.200 1.680 13.615 1.840 ;
        RECT  12.655 2.160 13.615 2.320 ;
        RECT  10.355 0.470 13.535 0.630 ;
        RECT  12.225 2.945 12.825 3.215 ;
        RECT  12.395 2.160 12.655 2.420 ;
        RECT  7.930 2.945 12.225 3.105 ;
        RECT  12.195 1.195 12.200 1.840 ;
        RECT  12.035 1.195 12.195 2.765 ;
        RECT  11.755 1.195 12.035 1.355 ;
        RECT  8.270 2.605 12.035 2.765 ;
        RECT  11.425 1.610 11.850 1.885 ;
        RECT  11.265 0.810 11.425 2.325 ;
        RECT  10.760 1.125 11.265 1.385 ;
        RECT  11.250 2.165 11.265 2.325 ;
        RECT  10.990 2.165 11.250 2.425 ;
        RECT  10.370 1.650 11.080 1.910 ;
        RECT  9.905 2.265 10.990 2.425 ;
        RECT  10.370 0.925 10.415 1.085 ;
        RECT  10.210 0.925 10.370 1.995 ;
        RECT  10.195 0.470 10.355 0.745 ;
        RECT  10.155 0.925 10.210 1.085 ;
        RECT  9.430 1.835 10.210 1.995 ;
        RECT  9.585 0.585 10.195 0.745 ;
        RECT  9.645 2.210 9.905 2.425 ;
        RECT  9.425 0.585 9.585 1.100 ;
        RECT  9.170 1.735 9.430 1.995 ;
        RECT  8.710 0.940 9.425 1.100 ;
        RECT  9.085 0.500 9.245 0.760 ;
        RECT  8.270 0.600 9.085 0.760 ;
        RECT  8.450 0.940 8.710 1.245 ;
        RECT  8.110 0.600 8.270 2.765 ;
        RECT  7.770 0.495 7.930 3.105 ;
        RECT  7.625 0.495 7.770 0.755 ;
        RECT  6.450 2.945 7.770 3.105 ;
        RECT  7.575 1.005 7.590 2.155 ;
        RECT  7.455 1.005 7.575 2.190 ;
        RECT  7.430 1.005 7.455 2.740 ;
        RECT  7.315 1.005 7.430 1.265 ;
        RECT  7.295 1.895 7.430 2.740 ;
        RECT  7.145 2.580 7.295 2.740 ;
        RECT  7.110 1.450 7.250 1.710 ;
        RECT  6.950 0.995 7.110 2.225 ;
        RECT  6.510 0.995 6.950 1.155 ;
        RECT  6.775 2.065 6.950 2.225 ;
        RECT  6.615 2.065 6.775 2.325 ;
        RECT  6.250 0.895 6.510 1.155 ;
        RECT  6.290 2.510 6.450 3.105 ;
        RECT  5.080 2.510 6.290 2.670 ;
        RECT  4.700 2.860 5.670 3.020 ;
        RECT  5.460 2.170 5.530 2.330 ;
        RECT  5.270 2.075 5.460 2.330 ;
        RECT  4.965 2.075 5.270 2.235 ;
        RECT  4.965 1.045 5.185 1.305 ;
        RECT  4.920 2.415 5.080 2.670 ;
        RECT  4.925 1.045 4.965 2.235 ;
        RECT  4.805 1.145 4.925 2.235 ;
        RECT  3.580 2.415 4.920 2.575 ;
        RECT  4.460 1.635 4.805 1.895 ;
        RECT  4.540 2.755 4.700 3.020 ;
        RECT  4.075 1.025 4.625 1.285 ;
        RECT  3.920 2.755 4.540 2.915 ;
        RECT  4.075 2.075 4.520 2.235 ;
        RECT  3.915 0.810 4.075 2.235 ;
        RECT  3.760 2.755 3.920 3.220 ;
        RECT  1.815 0.810 3.915 0.970 ;
        RECT  1.250 3.060 3.760 3.220 ;
        RECT  3.580 1.155 3.735 1.315 ;
        RECT  3.420 1.155 3.580 2.820 ;
        RECT  1.730 2.660 3.420 2.820 ;
        RECT  2.985 1.250 3.145 2.480 ;
        RECT  2.240 2.220 2.985 2.380 ;
        RECT  2.240 1.250 2.245 1.510 ;
        RECT  2.080 1.250 2.240 2.480 ;
        RECT  1.985 1.250 2.080 1.510 ;
        RECT  1.980 2.220 2.080 2.480 ;
        RECT  1.730 1.170 1.735 1.430 ;
        RECT  1.570 1.170 1.730 2.820 ;
        RECT  1.475 1.170 1.570 1.430 ;
        RECT  1.470 2.420 1.570 2.680 ;
        RECT  1.090 2.580 1.250 3.220 ;
        RECT  0.385 2.580 1.090 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.520 ;
    END
END SEDFFHQX8

MACRO SEDFFHQX4
    CLASS CORE ;
    FOREIGN SEDFFHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.700 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.990 1.255 2.400 ;
        RECT  0.975 1.565 1.235 2.400 ;
        END
        ANTENNAGATEAREA     0.1417 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.335 6.305 1.495 ;
        RECT  5.740 1.105 5.855 1.495 ;
        RECT  5.580 0.650 5.740 1.495 ;
        RECT  4.415 0.650 5.580 0.810 ;
        RECT  4.255 0.470 4.415 0.810 ;
        RECT  1.505 0.470 4.255 0.630 ;
        RECT  1.435 0.430 1.505 0.630 ;
        RECT  1.230 0.430 1.435 0.745 ;
        RECT  0.795 0.585 1.230 0.745 ;
        RECT  0.715 0.585 0.795 1.680 ;
        RECT  0.635 0.585 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1625 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.930 1.515 20.115 1.765 ;
        RECT  19.670 0.695 19.930 2.920 ;
        RECT  19.595 1.695 19.670 2.400 ;
        RECT  19.445 1.700 19.595 2.400 ;
        END
        ANTENNADIFFAREA     0.7980 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.855 1.725 6.770 1.885 ;
        RECT  5.645 1.700 5.855 1.990 ;
        RECT  5.335 1.700 5.645 1.860 ;
        RECT  5.175 1.575 5.335 1.860 ;
        END
        ANTENNAGATEAREA     0.1235 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.670 2.805 2.030 ;
        END
        ANTENNAGATEAREA     0.2834 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 1.290 9.995 1.580 ;
        RECT  9.815 1.155 9.975 1.580 ;
        RECT  9.585 1.290 9.815 1.580 ;
        END
        ANTENNAGATEAREA     0.4160 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.440 -0.250 20.700 0.250 ;
        RECT  20.180 -0.250 20.440 1.115 ;
        RECT  19.415 -0.250 20.180 0.250 ;
        RECT  19.155 -0.250 19.415 1.295 ;
        RECT  18.630 -0.250 19.155 0.250 ;
        RECT  18.370 -0.250 18.630 0.405 ;
        RECT  9.835 -0.250 18.370 0.250 ;
        RECT  9.575 -0.250 9.835 0.405 ;
        RECT  8.785 -0.250 9.575 0.250 ;
        RECT  8.525 -0.250 8.785 0.405 ;
        RECT  7.095 -0.250 8.525 0.250 ;
        RECT  6.835 -0.250 7.095 0.405 ;
        RECT  6.075 -0.250 6.835 0.250 ;
        RECT  5.815 -0.250 6.075 0.405 ;
        RECT  4.855 -0.250 5.815 0.250 ;
        RECT  4.595 -0.250 4.855 0.405 ;
        RECT  0.815 -0.250 4.595 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.440 3.440 20.700 3.940 ;
        RECT  20.180 2.255 20.440 3.940 ;
        RECT  19.385 3.440 20.180 3.940 ;
        RECT  19.125 3.285 19.385 3.940 ;
        RECT  18.505 3.440 19.125 3.940 ;
        RECT  18.245 3.285 18.505 3.940 ;
        RECT  15.910 3.440 18.245 3.940 ;
        RECT  15.650 3.285 15.910 3.940 ;
        RECT  14.795 3.440 15.650 3.940 ;
        RECT  14.535 3.285 14.795 3.940 ;
        RECT  13.520 3.440 14.535 3.940 ;
        RECT  13.260 3.285 13.520 3.940 ;
        RECT  11.790 3.440 13.260 3.940 ;
        RECT  11.530 3.285 11.790 3.940 ;
        RECT  10.710 3.440 11.530 3.940 ;
        RECT  10.450 3.285 10.710 3.940 ;
        RECT  8.725 3.440 10.450 3.940 ;
        RECT  8.465 3.285 8.725 3.940 ;
        RECT  6.965 3.440 8.465 3.940 ;
        RECT  6.705 3.285 6.965 3.940 ;
        RECT  6.110 3.440 6.705 3.940 ;
        RECT  5.850 2.945 6.110 3.940 ;
        RECT  5.100 3.440 5.850 3.940 ;
        RECT  4.840 3.285 5.100 3.940 ;
        RECT  4.360 3.405 4.840 3.940 ;
        RECT  4.100 3.095 4.360 3.940 ;
        RECT  0.870 3.440 4.100 3.940 ;
        RECT  0.610 2.925 0.870 3.940 ;
        RECT  0.000 3.440 0.610 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.895 2.575 18.935 2.835 ;
        RECT  18.735 0.845 18.895 2.835 ;
        RECT  18.625 0.845 18.735 1.225 ;
        RECT  18.640 1.885 18.735 2.145 ;
        RECT  18.675 2.575 18.735 2.835 ;
        RECT  18.190 0.845 18.625 1.005 ;
        RECT  18.445 1.405 18.555 1.665 ;
        RECT  18.285 1.185 18.445 2.880 ;
        RECT  17.850 1.185 18.285 1.345 ;
        RECT  16.820 2.720 18.285 2.880 ;
        RECT  18.030 0.470 18.190 1.005 ;
        RECT  17.945 1.530 18.105 2.535 ;
        RECT  14.490 0.470 18.030 0.630 ;
        RECT  17.510 1.530 17.945 1.690 ;
        RECT  17.360 2.375 17.945 2.535 ;
        RECT  17.690 0.910 17.850 1.345 ;
        RECT  17.605 1.875 17.765 2.190 ;
        RECT  17.360 0.910 17.690 1.070 ;
        RECT  17.170 1.875 17.605 2.035 ;
        RECT  17.335 3.060 17.595 3.260 ;
        RECT  17.350 1.250 17.510 1.690 ;
        RECT  17.100 0.810 17.360 1.070 ;
        RECT  17.200 2.220 17.360 2.535 ;
        RECT  16.820 1.250 17.350 1.410 ;
        RECT  16.250 3.060 17.335 3.220 ;
        RECT  16.820 2.220 17.200 2.380 ;
        RECT  17.010 1.635 17.170 2.035 ;
        RECT  16.230 0.810 17.100 0.970 ;
        RECT  15.540 1.635 17.010 1.795 ;
        RECT  16.560 1.155 16.820 1.410 ;
        RECT  16.560 2.120 16.820 2.380 ;
        RECT  16.660 2.565 16.820 2.880 ;
        RECT  16.280 2.565 16.660 2.725 ;
        RECT  15.880 1.250 16.560 1.410 ;
        RECT  15.370 2.120 16.560 2.280 ;
        RECT  16.020 2.465 16.280 2.725 ;
        RECT  16.090 2.940 16.250 3.220 ;
        RECT  16.070 0.810 16.230 1.070 ;
        RECT  14.160 2.940 16.090 3.100 ;
        RECT  15.720 0.910 15.880 1.410 ;
        RECT  15.370 0.910 15.720 1.070 ;
        RECT  15.380 1.250 15.540 1.795 ;
        RECT  14.760 1.250 15.380 1.410 ;
        RECT  15.110 0.810 15.370 1.070 ;
        RECT  15.110 2.120 15.370 2.760 ;
        RECT  14.940 1.635 15.200 1.850 ;
        RECT  14.340 2.600 15.110 2.760 ;
        RECT  13.955 1.690 14.940 1.850 ;
        RECT  14.600 0.810 14.760 1.410 ;
        RECT  14.145 0.810 14.600 0.970 ;
        RECT  14.330 0.430 14.490 0.630 ;
        RECT  13.695 0.430 14.330 0.590 ;
        RECT  14.000 2.605 14.160 3.100 ;
        RECT  13.885 0.770 14.145 0.970 ;
        RECT  12.195 2.605 14.000 2.765 ;
        RECT  13.875 1.150 13.955 2.320 ;
        RECT  11.425 0.810 13.885 0.970 ;
        RECT  13.795 1.150 13.875 2.425 ;
        RECT  12.435 1.150 13.795 1.310 ;
        RECT  13.615 2.160 13.795 2.425 ;
        RECT  13.535 0.430 13.695 0.630 ;
        RECT  12.200 1.680 13.615 1.840 ;
        RECT  12.655 2.160 13.615 2.320 ;
        RECT  10.355 0.470 13.535 0.630 ;
        RECT  12.225 2.945 12.825 3.215 ;
        RECT  12.395 2.160 12.655 2.420 ;
        RECT  7.930 2.945 12.225 3.105 ;
        RECT  12.195 1.195 12.200 1.840 ;
        RECT  12.035 1.195 12.195 2.765 ;
        RECT  11.755 1.195 12.035 1.355 ;
        RECT  8.270 2.605 12.035 2.765 ;
        RECT  11.425 1.610 11.850 1.885 ;
        RECT  11.265 0.810 11.425 2.325 ;
        RECT  10.760 1.125 11.265 1.385 ;
        RECT  11.250 2.165 11.265 2.325 ;
        RECT  10.990 2.165 11.250 2.425 ;
        RECT  10.370 1.650 11.080 1.910 ;
        RECT  9.905 2.265 10.990 2.425 ;
        RECT  10.370 0.925 10.415 1.085 ;
        RECT  10.210 0.925 10.370 1.995 ;
        RECT  10.195 0.470 10.355 0.745 ;
        RECT  10.155 0.925 10.210 1.085 ;
        RECT  9.430 1.835 10.210 1.995 ;
        RECT  9.585 0.585 10.195 0.745 ;
        RECT  9.645 2.210 9.905 2.425 ;
        RECT  9.425 0.585 9.585 1.100 ;
        RECT  9.170 1.735 9.430 1.995 ;
        RECT  8.710 0.940 9.425 1.100 ;
        RECT  9.085 0.500 9.245 0.760 ;
        RECT  8.270 0.600 9.085 0.760 ;
        RECT  8.450 0.940 8.710 1.245 ;
        RECT  8.110 0.600 8.270 2.765 ;
        RECT  7.770 0.495 7.930 3.105 ;
        RECT  7.625 0.495 7.770 0.755 ;
        RECT  6.450 2.945 7.770 3.105 ;
        RECT  7.575 1.005 7.590 2.155 ;
        RECT  7.455 1.005 7.575 2.190 ;
        RECT  7.430 1.005 7.455 2.740 ;
        RECT  7.315 1.005 7.430 1.265 ;
        RECT  7.295 1.895 7.430 2.740 ;
        RECT  7.145 2.580 7.295 2.740 ;
        RECT  7.110 1.450 7.250 1.710 ;
        RECT  6.950 0.995 7.110 2.225 ;
        RECT  6.510 0.995 6.950 1.155 ;
        RECT  6.775 2.065 6.950 2.225 ;
        RECT  6.615 2.065 6.775 2.325 ;
        RECT  6.250 0.895 6.510 1.155 ;
        RECT  6.290 2.510 6.450 3.105 ;
        RECT  5.080 2.510 6.290 2.670 ;
        RECT  4.700 2.860 5.670 3.020 ;
        RECT  5.460 2.170 5.530 2.330 ;
        RECT  5.270 2.075 5.460 2.330 ;
        RECT  4.965 2.075 5.270 2.235 ;
        RECT  4.965 1.045 5.185 1.305 ;
        RECT  4.920 2.415 5.080 2.670 ;
        RECT  4.925 1.045 4.965 2.235 ;
        RECT  4.805 1.145 4.925 2.235 ;
        RECT  3.580 2.415 4.920 2.575 ;
        RECT  4.460 1.635 4.805 1.895 ;
        RECT  4.540 2.755 4.700 3.020 ;
        RECT  4.075 1.025 4.625 1.285 ;
        RECT  3.920 2.755 4.540 2.915 ;
        RECT  4.075 2.075 4.520 2.235 ;
        RECT  3.915 0.810 4.075 2.235 ;
        RECT  3.760 2.755 3.920 3.220 ;
        RECT  1.815 0.810 3.915 0.970 ;
        RECT  1.250 3.060 3.760 3.220 ;
        RECT  3.580 1.155 3.735 1.315 ;
        RECT  3.420 1.155 3.580 2.820 ;
        RECT  1.730 2.660 3.420 2.820 ;
        RECT  2.985 1.250 3.145 2.480 ;
        RECT  2.240 2.220 2.985 2.380 ;
        RECT  2.240 1.250 2.245 1.510 ;
        RECT  2.080 1.250 2.240 2.480 ;
        RECT  1.985 1.250 2.080 1.510 ;
        RECT  1.980 2.220 2.080 2.480 ;
        RECT  1.730 1.170 1.735 1.430 ;
        RECT  1.570 1.170 1.730 2.820 ;
        RECT  1.475 1.170 1.570 1.430 ;
        RECT  1.470 2.420 1.570 2.680 ;
        RECT  1.090 2.580 1.250 3.220 ;
        RECT  0.385 2.580 1.090 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.255 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.520 ;
    END
END SEDFFHQX4

MACRO SEDFFHQX2
    CLASS CORE ;
    FOREIGN SEDFFHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.565 1.265 1.825 ;
        RECT  1.045 1.565 1.255 2.400 ;
        RECT  1.005 1.565 1.045 1.825 ;
        END
        ANTENNAGATEAREA     0.0754 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.890 1.335 5.255 1.495 ;
        RECT  4.730 1.000 4.890 1.495 ;
        RECT  4.450 1.000 4.730 1.160 ;
        RECT  4.290 0.620 4.450 1.160 ;
        RECT  2.955 0.620 4.290 0.780 ;
        RECT  2.795 0.490 2.955 0.780 ;
        RECT  2.455 0.490 2.795 0.650 ;
        RECT  2.295 0.430 2.455 0.650 ;
        RECT  1.670 0.430 2.295 0.590 ;
        RECT  1.510 0.430 1.670 0.735 ;
        RECT  1.505 0.575 1.510 0.735 ;
        RECT  1.230 0.575 1.505 0.835 ;
        RECT  0.795 0.675 1.230 0.835 ;
        RECT  0.715 0.675 0.795 1.680 ;
        RECT  0.635 0.675 0.715 1.730 ;
        RECT  0.585 1.105 0.635 1.730 ;
        RECT  0.455 1.470 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1378 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.860 1.105 15.975 2.585 ;
        RECT  15.820 1.105 15.860 2.895 ;
        RECT  15.660 0.695 15.820 2.895 ;
        RECT  15.560 0.695 15.660 1.295 ;
        RECT  15.600 1.955 15.660 2.895 ;
        RECT  15.305 2.520 15.600 2.810 ;
        END
        ANTENNADIFFAREA     0.7140 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.625 5.880 1.885 ;
        RECT  4.935 1.680 5.720 1.840 ;
        RECT  4.930 1.680 4.935 1.990 ;
        RECT  4.725 1.675 4.930 1.990 ;
        RECT  4.285 1.675 4.725 1.835 ;
        RECT  4.125 1.575 4.285 1.835 ;
        END
        ANTENNAGATEAREA     0.1001 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.535 2.635 1.990 ;
        RECT  2.305 1.535 2.425 1.895 ;
        END
        ANTENNAGATEAREA     0.1482 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 1.285 8.970 1.670 ;
        END
        ANTENNAGATEAREA     0.2327 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.270 -0.250 16.100 0.250 ;
        RECT  14.330 -0.250 15.270 0.405 ;
        RECT  9.010 -0.250 14.330 0.250 ;
        RECT  8.750 -0.250 9.010 0.405 ;
        RECT  7.710 -0.250 8.750 0.250 ;
        RECT  7.450 -0.250 7.710 0.405 ;
        RECT  6.370 -0.250 7.450 0.250 ;
        RECT  5.770 -0.250 6.370 0.405 ;
        RECT  4.880 -0.250 5.770 0.250 ;
        RECT  4.830 -0.250 4.880 0.405 ;
        RECT  4.670 -0.250 4.830 0.795 ;
        RECT  4.620 -0.250 4.670 0.405 ;
        RECT  3.395 -0.250 4.620 0.250 ;
        RECT  3.135 -0.250 3.395 0.405 ;
        RECT  0.815 -0.250 3.135 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.315 3.440 16.100 3.940 ;
        RECT  15.055 3.285 15.315 3.940 ;
        RECT  14.370 3.440 15.055 3.940 ;
        RECT  14.110 2.840 14.370 3.940 ;
        RECT  12.150 3.440 14.110 3.940 ;
        RECT  11.890 3.285 12.150 3.940 ;
        RECT  10.435 3.440 11.890 3.940 ;
        RECT  10.175 3.285 10.435 3.940 ;
        RECT  8.415 3.440 10.175 3.940 ;
        RECT  8.155 3.285 8.415 3.940 ;
        RECT  6.485 3.440 8.155 3.940 ;
        RECT  6.225 3.285 6.485 3.940 ;
        RECT  5.250 3.440 6.225 3.940 ;
        RECT  4.990 2.925 5.250 3.940 ;
        RECT  4.165 3.440 4.990 3.940 ;
        RECT  3.905 3.285 4.165 3.940 ;
        RECT  3.235 3.440 3.905 3.940 ;
        RECT  3.075 3.035 3.235 3.940 ;
        RECT  0.815 3.440 3.075 3.940 ;
        RECT  0.555 2.925 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.865 2.405 14.950 2.665 ;
        RECT  14.865 0.890 14.890 1.150 ;
        RECT  14.705 0.890 14.865 2.665 ;
        RECT  14.630 0.890 14.705 1.375 ;
        RECT  14.690 2.035 14.705 2.665 ;
        RECT  14.265 2.035 14.690 2.195 ;
        RECT  14.090 1.215 14.630 1.375 ;
        RECT  14.365 1.555 14.525 1.815 ;
        RECT  13.750 1.605 14.365 1.765 ;
        RECT  14.005 2.035 14.265 2.295 ;
        RECT  13.930 0.470 14.090 1.375 ;
        RECT  9.525 0.470 13.930 0.630 ;
        RECT  13.590 0.860 13.750 1.800 ;
        RECT  13.575 2.035 13.735 2.630 ;
        RECT  13.565 3.100 13.615 3.260 ;
        RECT  13.180 0.860 13.590 1.020 ;
        RECT  13.365 1.640 13.590 1.800 ;
        RECT  13.025 2.470 13.575 2.630 ;
        RECT  13.355 2.945 13.565 3.260 ;
        RECT  13.025 1.200 13.410 1.460 ;
        RECT  13.205 1.640 13.365 2.285 ;
        RECT  11.510 2.945 13.355 3.105 ;
        RECT  13.000 1.200 13.025 2.630 ;
        RECT  12.865 0.810 13.000 2.630 ;
        RECT  12.840 0.810 12.865 1.360 ;
        RECT  10.180 0.810 12.840 0.970 ;
        RECT  12.630 2.025 12.685 2.630 ;
        RECT  12.630 1.150 12.660 1.310 ;
        RECT  12.470 1.150 12.630 2.630 ;
        RECT  12.400 1.150 12.470 1.310 ;
        RECT  11.705 2.470 12.470 2.630 ;
        RECT  12.120 1.585 12.290 1.845 ;
        RECT  11.960 1.180 12.120 2.290 ;
        RECT  11.055 1.180 11.960 1.340 ;
        RECT  11.025 2.130 11.960 2.290 ;
        RECT  11.350 2.605 11.510 3.105 ;
        RECT  10.845 1.720 11.485 1.880 ;
        RECT  10.845 2.605 11.350 2.765 ;
        RECT  11.035 3.100 11.115 3.260 ;
        RECT  10.855 2.945 11.035 3.260 ;
        RECT  7.435 2.945 10.855 3.105 ;
        RECT  10.685 1.225 10.845 2.765 ;
        RECT  10.360 1.225 10.685 1.385 ;
        RECT  8.475 2.605 10.685 2.765 ;
        RECT  10.180 1.660 10.505 1.920 ;
        RECT  10.020 0.810 10.180 2.385 ;
        RECT  9.710 0.810 10.020 0.970 ;
        RECT  9.250 2.225 10.020 2.385 ;
        RECT  9.500 1.650 9.825 1.910 ;
        RECT  9.365 0.470 9.525 0.765 ;
        RECT  9.340 0.945 9.500 2.020 ;
        RECT  7.880 0.605 9.365 0.765 ;
        RECT  9.200 0.945 9.340 1.105 ;
        RECT  8.905 1.860 9.340 2.020 ;
        RECT  8.745 1.860 8.905 2.120 ;
        RECT  8.315 1.985 8.475 2.765 ;
        RECT  8.220 0.945 8.345 1.105 ;
        RECT  8.220 1.985 8.315 2.145 ;
        RECT  8.060 0.945 8.220 2.145 ;
        RECT  7.880 2.325 8.135 2.585 ;
        RECT  7.875 0.605 7.880 2.585 ;
        RECT  7.720 0.605 7.875 2.485 ;
        RECT  7.275 1.065 7.435 3.105 ;
        RECT  6.920 1.065 7.275 1.225 ;
        RECT  6.095 2.945 7.275 3.105 ;
        RECT  6.905 1.425 7.065 2.765 ;
        RECT  6.760 0.755 6.920 1.225 ;
        RECT  6.580 1.425 6.905 1.585 ;
        RECT  6.745 2.505 6.905 2.765 ;
        RECT  6.240 1.795 6.635 2.055 ;
        RECT  6.420 0.945 6.580 1.585 ;
        RECT  6.200 0.945 6.420 1.105 ;
        RECT  6.100 1.285 6.240 2.225 ;
        RECT  6.080 1.285 6.100 2.325 ;
        RECT  5.935 2.520 6.095 3.105 ;
        RECT  5.595 1.285 6.080 1.445 ;
        RECT  5.840 2.065 6.080 2.325 ;
        RECT  3.915 2.520 5.935 2.680 ;
        RECT  5.450 0.995 5.595 1.445 ;
        RECT  5.435 0.895 5.450 1.445 ;
        RECT  5.190 0.895 5.435 1.155 ;
        RECT  4.550 2.860 4.810 3.120 ;
        RECT  4.530 2.170 4.680 2.330 ;
        RECT  3.575 2.860 4.550 3.020 ;
        RECT  4.370 2.015 4.530 2.330 ;
        RECT  3.940 2.015 4.370 2.175 ;
        RECT  3.940 1.045 4.110 1.305 ;
        RECT  3.780 1.045 3.940 2.175 ;
        RECT  3.755 2.355 3.915 2.680 ;
        RECT  3.535 1.575 3.780 1.835 ;
        RECT  2.555 2.355 3.755 2.515 ;
        RECT  3.340 1.045 3.600 1.305 ;
        RECT  3.120 2.015 3.595 2.175 ;
        RECT  3.415 2.695 3.575 3.020 ;
        RECT  2.895 2.695 3.415 2.855 ;
        RECT  3.120 1.095 3.340 1.305 ;
        RECT  2.960 1.095 3.120 2.175 ;
        RECT  2.615 1.095 2.960 1.255 ;
        RECT  2.735 2.695 2.895 3.135 ;
        RECT  1.365 2.975 2.735 3.135 ;
        RECT  2.455 0.835 2.615 1.255 ;
        RECT  2.395 2.355 2.555 2.735 ;
        RECT  2.115 0.835 2.455 0.995 ;
        RECT  1.705 2.575 2.395 2.735 ;
        RECT  2.115 1.175 2.275 1.335 ;
        RECT  2.115 2.130 2.215 2.390 ;
        RECT  1.850 0.770 2.115 0.995 ;
        RECT  1.955 1.175 2.115 2.390 ;
        RECT  1.705 1.210 1.725 1.470 ;
        RECT  1.545 1.210 1.705 2.735 ;
        RECT  1.515 1.210 1.545 2.390 ;
        RECT  1.465 1.210 1.515 1.470 ;
        RECT  1.445 2.130 1.515 2.390 ;
        RECT  1.205 2.580 1.365 3.135 ;
        RECT  0.385 2.580 1.205 2.740 ;
        RECT  0.275 1.025 0.385 1.285 ;
        RECT  0.275 2.185 0.385 2.740 ;
        RECT  0.225 1.025 0.275 2.740 ;
        RECT  0.115 1.025 0.225 2.450 ;
    END
END SEDFFHQX2

MACRO SEDFFHQX1
    CLASS CORE ;
    FOREIGN SEDFFHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 1.925 1.255 2.400 ;
        RECT  1.055 1.565 1.215 2.400 ;
        RECT  1.045 1.925 1.055 2.400 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.455 4.885 1.615 ;
        RECT  4.420 0.745 4.580 1.615 ;
        RECT  4.265 0.745 4.420 1.355 ;
        RECT  2.975 0.745 4.265 0.905 ;
        RECT  2.815 0.470 2.975 0.905 ;
        RECT  1.530 0.470 2.815 0.630 ;
        RECT  1.230 0.470 1.530 0.805 ;
        RECT  0.795 0.645 1.230 0.805 ;
        RECT  0.665 0.645 0.795 1.580 ;
        RECT  0.610 0.645 0.665 1.730 ;
        RECT  0.585 1.105 0.610 1.730 ;
        RECT  0.505 1.355 0.585 1.730 ;
        END
        ANTENNAGATEAREA     0.1274 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.540 1.515 14.595 2.585 ;
        RECT  14.395 1.060 14.540 2.810 ;
        RECT  14.380 1.010 14.395 2.810 ;
        RECT  14.235 1.010 14.380 1.270 ;
        RECT  14.220 2.525 14.380 2.810 ;
        RECT  14.135 2.525 14.220 3.170 ;
        RECT  13.960 2.520 14.135 3.170 ;
        RECT  13.925 2.520 13.960 2.995 ;
        END
        ANTENNADIFFAREA     0.5262 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.155 1.675 5.315 1.955 ;
        RECT  4.015 1.795 5.155 1.955 ;
        RECT  3.805 1.700 4.015 2.010 ;
        END
        ANTENNAGATEAREA     0.0975 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.520 2.635 1.990 ;
        RECT  2.295 1.520 2.425 1.920 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.290 7.695 1.905 ;
        END
        ANTENNAGATEAREA     0.1430 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.580 -0.250 14.720 0.250 ;
        RECT  13.320 -0.250 13.580 0.405 ;
        RECT  9.465 -0.250 13.320 0.250 ;
        RECT  9.205 -0.250 9.465 0.405 ;
        RECT  8.575 -0.250 9.205 0.250 ;
        RECT  8.315 -0.250 8.575 0.405 ;
        RECT  7.135 -0.250 8.315 0.250 ;
        RECT  6.875 -0.250 7.135 0.405 ;
        RECT  5.580 -0.250 6.875 0.250 ;
        RECT  5.320 -0.250 5.580 0.405 ;
        RECT  4.715 -0.250 5.320 0.250 ;
        RECT  4.455 -0.250 4.715 0.405 ;
        RECT  3.440 -0.250 4.455 0.250 ;
        RECT  3.180 -0.250 3.440 0.405 ;
        RECT  0.815 -0.250 3.180 0.250 ;
        RECT  0.555 -0.250 0.815 0.405 ;
        RECT  0.000 -0.250 0.555 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.620 3.440 14.720 3.940 ;
        RECT  13.360 2.610 13.620 3.940 ;
        RECT  11.645 3.440 13.360 3.940 ;
        RECT  11.385 3.285 11.645 3.940 ;
        RECT  6.945 3.440 11.385 3.940 ;
        RECT  6.685 3.285 6.945 3.940 ;
        RECT  4.825 3.440 6.685 3.940 ;
        RECT  4.565 2.945 4.825 3.940 ;
        RECT  3.815 3.440 4.565 3.940 ;
        RECT  3.555 2.945 3.815 3.940 ;
        RECT  2.575 3.440 3.555 3.940 ;
        RECT  2.315 2.780 2.575 3.940 ;
        RECT  0.815 3.440 2.315 3.940 ;
        RECT  0.555 3.285 0.815 3.940 ;
        RECT  0.000 3.440 0.555 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.055 2.000 14.200 2.260 ;
        RECT  14.055 0.430 14.175 0.590 ;
        RECT  14.040 0.430 14.055 2.260 ;
        RECT  13.895 0.430 14.040 2.160 ;
        RECT  12.785 0.585 13.895 0.745 ;
        RECT  13.400 2.000 13.895 2.160 ;
        RECT  13.550 1.380 13.710 1.645 ;
        RECT  13.370 1.380 13.550 1.540 ;
        RECT  13.240 1.895 13.400 2.160 ;
        RECT  13.210 0.925 13.370 1.540 ;
        RECT  12.535 0.925 13.210 1.085 ;
        RECT  12.995 2.975 13.080 3.235 ;
        RECT  12.835 1.265 12.995 3.235 ;
        RECT  12.760 1.265 12.835 1.525 ;
        RECT  12.820 2.915 12.835 3.235 ;
        RECT  10.855 2.915 12.820 3.075 ;
        RECT  12.625 0.470 12.785 0.745 ;
        RECT  12.535 2.410 12.655 2.670 ;
        RECT  9.805 0.470 12.625 0.630 ;
        RECT  12.375 0.925 12.535 2.670 ;
        RECT  12.360 1.130 12.375 1.390 ;
        RECT  12.090 2.475 12.195 2.735 ;
        RECT  10.150 0.810 12.180 0.970 ;
        RECT  11.930 1.195 12.090 2.735 ;
        RECT  11.660 1.195 11.930 1.355 ;
        RECT  11.165 2.575 11.930 2.735 ;
        RECT  11.235 1.845 11.750 2.105 ;
        RECT  11.075 1.185 11.235 2.395 ;
        RECT  10.330 1.185 11.075 1.345 ;
        RECT  10.695 2.235 11.075 2.395 ;
        RECT  10.355 1.890 10.895 2.050 ;
        RECT  10.695 2.720 10.855 3.075 ;
        RECT  10.535 2.235 10.695 2.540 ;
        RECT  10.355 2.720 10.695 2.880 ;
        RECT  7.285 3.060 10.515 3.220 ;
        RECT  10.195 1.545 10.355 2.880 ;
        RECT  9.760 1.545 10.195 1.705 ;
        RECT  7.625 2.720 10.195 2.880 ;
        RECT  9.990 0.810 10.150 1.150 ;
        RECT  9.390 1.895 10.015 2.055 ;
        RECT  9.390 0.990 9.990 1.150 ;
        RECT  9.645 0.470 9.805 0.760 ;
        RECT  9.600 1.365 9.760 1.705 ;
        RECT  6.875 0.600 9.645 0.760 ;
        RECT  9.230 0.990 9.390 2.540 ;
        RECT  8.850 0.990 9.230 1.250 ;
        RECT  7.965 2.380 9.230 2.540 ;
        RECT  8.420 1.500 9.050 1.760 ;
        RECT  8.260 1.135 8.420 2.165 ;
        RECT  8.140 1.135 8.260 1.295 ;
        RECT  8.160 2.005 8.260 2.165 ;
        RECT  7.880 1.035 8.140 1.295 ;
        RECT  7.805 2.125 7.965 2.540 ;
        RECT  7.465 2.605 7.625 2.880 ;
        RECT  7.265 0.950 7.610 1.110 ;
        RECT  7.265 2.605 7.465 2.765 ;
        RECT  7.125 2.945 7.285 3.220 ;
        RECT  7.105 0.950 7.265 2.765 ;
        RECT  6.505 2.945 7.125 3.105 ;
        RECT  6.715 0.600 6.875 1.720 ;
        RECT  6.505 2.150 6.535 2.410 ;
        RECT  6.345 0.720 6.505 3.220 ;
        RECT  6.245 0.720 6.345 0.880 ;
        RECT  5.165 3.060 6.345 3.220 ;
        RECT  5.985 0.620 6.245 0.880 ;
        RECT  6.005 1.180 6.165 2.875 ;
        RECT  5.900 1.180 6.005 1.340 ;
        RECT  5.735 2.715 6.005 2.875 ;
        RECT  5.655 1.500 5.795 1.760 ;
        RECT  5.495 1.085 5.655 2.295 ;
        RECT  4.890 1.085 5.495 1.245 ;
        RECT  5.275 2.135 5.495 2.295 ;
        RECT  5.005 2.605 5.165 3.220 ;
        RECT  2.915 2.605 5.005 2.765 ;
        RECT  3.605 2.240 4.245 2.400 ;
        RECT  3.605 1.085 3.815 1.245 ;
        RECT  3.445 1.085 3.605 2.400 ;
        RECT  3.155 1.590 3.445 1.850 ;
        RECT  2.975 1.130 3.255 1.390 ;
        RECT  2.975 2.100 3.255 2.260 ;
        RECT  2.815 1.130 2.975 2.260 ;
        RECT  2.755 2.440 2.915 2.765 ;
        RECT  2.635 1.130 2.815 1.290 ;
        RECT  1.655 2.440 2.755 2.600 ;
        RECT  2.475 0.810 2.635 1.290 ;
        RECT  1.835 0.810 2.475 0.970 ;
        RECT  2.115 1.180 2.295 1.340 ;
        RECT  2.115 2.100 2.215 2.260 ;
        RECT  1.955 1.180 2.115 2.260 ;
        RECT  1.505 2.780 1.765 3.035 ;
        RECT  1.495 1.130 1.655 2.600 ;
        RECT  0.385 2.780 1.505 2.940 ;
        RECT  0.325 2.255 0.385 2.940 ;
        RECT  0.325 1.025 0.335 1.285 ;
        RECT  0.225 1.025 0.325 2.940 ;
        RECT  0.165 1.025 0.225 2.515 ;
        RECT  0.125 2.255 0.165 2.515 ;
    END
END SEDFFHQX1

MACRO SDFFSRHQX8
    CLASS CORE ;
    FOREIGN SDFFSRHQX8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.320 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.655 7.695 2.400 ;
        RECT  7.435 1.655 7.485 1.915 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.185 1.265 6.375 2.080 ;
        RECT  5.965 1.265 6.185 1.635 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 1.615 5.445 1.875 ;
        RECT  5.180 1.615 5.340 2.540 ;
        RECT  2.755 2.380 5.180 2.540 ;
        RECT  2.595 1.620 2.755 2.540 ;
        RECT  2.425 1.700 2.595 2.175 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.165 1.525 14.425 1.785 ;
        RECT  13.215 1.625 14.165 1.785 ;
        RECT  12.845 1.625 13.215 1.990 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.735 0.980 19.195 2.395 ;
        RECT  18.685 0.980 18.735 2.585 ;
        RECT  18.525 0.690 18.685 3.045 ;
        RECT  18.425 0.690 18.525 1.290 ;
        RECT  18.425 1.990 18.525 3.045 ;
        RECT  17.665 0.980 18.425 1.290 ;
        RECT  18.275 1.990 18.425 2.400 ;
        RECT  17.665 1.990 18.275 2.395 ;
        RECT  17.405 0.690 17.665 1.290 ;
        RECT  17.405 1.990 17.665 3.045 ;
        END
        ANTENNADIFFAREA     1.6264 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.290 4.265 1.580 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.335 2.185 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 -0.250 19.320 0.250 ;
        RECT  18.935 -0.250 19.195 0.755 ;
        RECT  18.175 -0.250 18.935 0.250 ;
        RECT  17.915 -0.250 18.175 0.755 ;
        RECT  17.125 -0.250 17.915 0.250 ;
        RECT  16.865 -0.250 17.125 1.135 ;
        RECT  16.525 -0.250 16.865 0.405 ;
        RECT  15.115 -0.250 16.525 0.250 ;
        RECT  14.855 -0.250 15.115 0.405 ;
        RECT  12.070 -0.250 14.855 0.250 ;
        RECT  11.810 -0.250 12.070 0.405 ;
        RECT  9.830 -0.250 11.810 0.250 ;
        RECT  9.230 -0.250 9.830 0.405 ;
        RECT  7.615 -0.250 9.230 0.250 ;
        RECT  7.355 -0.250 7.615 0.405 ;
        RECT  6.595 -0.250 7.355 0.250 ;
        RECT  5.995 -0.250 6.595 0.405 ;
        RECT  4.115 -0.250 5.995 0.250 ;
        RECT  3.875 -0.250 4.115 0.405 ;
        RECT  3.515 -0.250 3.875 0.745 ;
        RECT  0.940 -0.250 3.515 0.250 ;
        RECT  0.340 -0.250 0.940 0.405 ;
        RECT  0.000 -0.250 0.340 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 3.440 19.320 3.940 ;
        RECT  18.935 2.615 19.195 3.940 ;
        RECT  18.175 3.440 18.935 3.940 ;
        RECT  17.915 2.615 18.175 3.940 ;
        RECT  17.155 3.440 17.915 3.940 ;
        RECT  16.895 2.275 17.155 3.940 ;
        RECT  16.215 2.955 16.895 3.940 ;
        RECT  14.775 3.440 16.215 3.940 ;
        RECT  14.515 3.285 14.775 3.940 ;
        RECT  12.135 3.440 14.515 3.940 ;
        RECT  11.875 3.285 12.135 3.940 ;
        RECT  10.990 3.440 11.875 3.940 ;
        RECT  10.730 3.285 10.990 3.940 ;
        RECT  9.460 3.440 10.730 3.940 ;
        RECT  9.200 2.660 9.460 3.940 ;
        RECT  6.920 3.440 9.200 3.940 ;
        RECT  6.660 3.285 6.920 3.940 ;
        RECT  1.380 3.440 6.660 3.940 ;
        RECT  0.780 3.285 1.380 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.325 1.510 18.055 1.770 ;
        RECT  16.665 1.495 17.325 1.770 ;
        RECT  16.505 0.680 16.665 2.580 ;
        RECT  15.655 0.680 16.505 0.840 ;
        RECT  16.435 1.510 16.505 1.770 ;
        RECT  15.725 2.420 16.505 2.580 ;
        RECT  16.225 1.035 16.325 1.295 ;
        RECT  16.225 1.955 16.325 2.215 ;
        RECT  16.065 1.035 16.225 2.215 ;
        RECT  15.695 1.725 16.065 1.985 ;
        RECT  15.565 2.420 15.725 2.935 ;
        RECT  15.495 0.680 15.655 1.025 ;
        RECT  13.825 2.775 15.565 2.935 ;
        RECT  15.395 0.765 15.495 1.025 ;
        RECT  15.385 1.205 15.485 1.465 ;
        RECT  13.315 0.840 15.395 1.000 ;
        RECT  15.285 1.205 15.385 2.295 ;
        RECT  15.225 1.205 15.285 2.595 ;
        RECT  15.125 2.035 15.225 2.595 ;
        RECT  14.115 2.435 15.125 2.595 ;
        RECT  14.805 1.995 14.905 2.255 ;
        RECT  14.645 1.180 14.805 2.255 ;
        RECT  13.095 1.180 14.645 1.340 ;
        RECT  13.955 2.055 14.115 2.595 ;
        RECT  13.825 2.055 13.955 2.330 ;
        RECT  13.095 0.470 13.945 0.630 ;
        RECT  12.665 2.170 13.825 2.330 ;
        RECT  13.565 2.775 13.825 3.035 ;
        RECT  12.660 2.510 13.260 2.770 ;
        RECT  12.935 0.470 13.095 1.340 ;
        RECT  12.475 3.060 13.055 3.220 ;
        RECT  12.415 0.470 12.935 0.630 ;
        RECT  12.665 0.810 12.755 1.085 ;
        RECT  12.595 0.810 12.665 2.330 ;
        RECT  11.585 2.510 12.660 2.670 ;
        RECT  12.505 0.925 12.595 2.330 ;
        RECT  11.290 0.925 12.505 1.085 ;
        RECT  12.005 2.015 12.505 2.330 ;
        RECT  12.315 2.945 12.475 3.220 ;
        RECT  12.255 0.470 12.415 0.745 ;
        RECT  12.155 1.265 12.315 1.525 ;
        RECT  10.450 2.945 12.315 3.105 ;
        RECT  11.630 0.585 12.255 0.745 ;
        RECT  10.950 1.265 12.155 1.425 ;
        RECT  11.470 0.470 11.630 0.745 ;
        RECT  11.325 2.460 11.585 2.720 ;
        RECT  10.170 0.470 11.470 0.630 ;
        RECT  10.960 2.460 11.325 2.620 ;
        RECT  11.130 0.810 11.290 1.085 ;
        RECT  10.510 0.810 11.130 0.970 ;
        RECT  10.950 1.920 10.960 2.620 ;
        RECT  10.800 1.150 10.950 2.620 ;
        RECT  10.790 1.150 10.800 2.130 ;
        RECT  10.690 1.150 10.790 1.425 ;
        RECT  10.675 1.870 10.790 2.130 ;
        RECT  10.350 0.810 10.510 1.145 ;
        RECT  10.350 1.385 10.510 1.645 ;
        RECT  10.190 2.945 10.450 3.245 ;
        RECT  7.250 0.985 10.350 1.145 ;
        RECT  10.230 1.485 10.350 1.645 ;
        RECT  10.230 2.390 10.280 2.650 ;
        RECT  10.070 1.485 10.230 2.650 ;
        RECT  9.800 2.945 10.190 3.105 ;
        RECT  10.010 0.470 10.170 0.745 ;
        RECT  9.075 1.485 10.070 1.645 ;
        RECT  10.020 2.390 10.070 2.650 ;
        RECT  9.335 0.585 10.010 0.745 ;
        RECT  9.640 2.210 9.800 3.105 ;
        RECT  8.720 2.210 9.640 2.370 ;
        RECT  9.075 0.585 9.335 0.805 ;
        RECT  4.215 0.585 9.075 0.745 ;
        RECT  8.815 1.325 9.075 1.645 ;
        RECT  8.035 1.485 8.815 1.645 ;
        RECT  8.560 1.925 8.720 3.220 ;
        RECT  8.375 1.925 8.560 2.085 ;
        RECT  7.260 3.060 8.560 3.220 ;
        RECT  7.600 2.720 8.380 2.880 ;
        RECT  8.215 1.825 8.375 2.085 ;
        RECT  8.035 2.350 8.240 2.510 ;
        RECT  7.875 1.485 8.035 2.510 ;
        RECT  7.440 2.605 7.600 2.880 ;
        RECT  6.715 2.605 7.440 2.765 ;
        RECT  7.250 2.265 7.290 2.425 ;
        RECT  7.100 2.945 7.260 3.220 ;
        RECT  7.090 0.935 7.250 2.425 ;
        RECT  6.480 2.945 7.100 3.105 ;
        RECT  6.895 0.935 7.090 1.195 ;
        RECT  7.030 2.265 7.090 2.425 ;
        RECT  6.555 0.925 6.715 2.765 ;
        RECT  5.215 0.925 6.555 1.085 ;
        RECT  5.860 2.395 6.555 2.655 ;
        RECT  6.320 2.945 6.480 3.220 ;
        RECT  1.725 3.060 6.320 3.220 ;
        RECT  5.785 1.865 6.005 2.215 ;
        RECT  5.680 1.275 5.785 2.215 ;
        RECT  5.625 1.275 5.680 2.880 ;
        RECT  4.965 1.275 5.625 1.435 ;
        RECT  5.520 2.055 5.625 2.880 ;
        RECT  2.235 2.720 5.520 2.880 ;
        RECT  4.955 0.925 5.215 1.095 ;
        RECT  4.605 2.040 5.000 2.200 ;
        RECT  4.785 1.275 4.965 1.560 ;
        RECT  4.605 0.925 4.655 1.085 ;
        RECT  4.445 0.925 4.605 2.200 ;
        RECT  4.395 0.925 4.445 1.085 ;
        RECT  4.055 0.585 4.215 1.110 ;
        RECT  3.235 0.950 4.055 1.110 ;
        RECT  3.235 2.040 4.050 2.200 ;
        RECT  3.075 0.930 3.235 2.200 ;
        RECT  2.975 0.930 3.075 1.190 ;
        RECT  2.765 0.470 2.975 0.750 ;
        RECT  2.575 0.930 2.975 1.090 ;
        RECT  1.285 0.470 2.765 0.630 ;
        RECT  2.415 0.810 2.575 1.090 ;
        RECT  1.625 0.810 2.415 0.970 ;
        RECT  2.075 1.150 2.235 2.880 ;
        RECT  1.805 1.150 2.075 1.310 ;
        RECT  1.625 1.575 1.895 1.835 ;
        RECT  1.565 2.120 1.725 3.220 ;
        RECT  1.465 0.810 1.625 1.835 ;
        RECT  1.465 2.120 1.565 2.380 ;
        RECT  1.295 1.575 1.465 1.835 ;
        RECT  1.015 2.120 1.465 2.280 ;
        RECT  1.125 0.470 1.285 0.745 ;
        RECT  1.125 0.970 1.285 1.230 ;
        RECT  0.675 0.585 1.125 0.745 ;
        RECT  1.015 1.070 1.125 1.230 ;
        RECT  0.855 1.070 1.015 2.280 ;
        RECT  0.515 0.585 0.675 2.895 ;
        RECT  0.125 0.835 0.515 1.095 ;
        RECT  0.385 2.735 0.515 2.895 ;
        RECT  0.125 2.735 0.385 2.995 ;
    END
END SDFFSRHQX8

MACRO SDFFSRHQX4
    CLASS CORE ;
    FOREIGN SDFFSRHQX4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.940 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 1.655 7.695 2.400 ;
        RECT  7.435 1.655 7.485 1.915 ;
        END
        ANTENNAGATEAREA     0.2691 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.185 1.265 6.375 2.080 ;
        RECT  5.965 1.265 6.185 1.635 ;
        END
        ANTENNAGATEAREA     0.1547 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.340 1.615 5.445 1.875 ;
        RECT  5.180 1.615 5.340 2.540 ;
        RECT  2.755 2.380 5.180 2.540 ;
        RECT  2.595 1.620 2.755 2.540 ;
        RECT  2.425 1.700 2.595 2.175 ;
        END
        ANTENNAGATEAREA     0.2600 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.295 1.525 14.455 1.820 ;
        RECT  13.215 1.660 14.295 1.820 ;
        RECT  13.125 1.660 13.215 1.990 ;
        RECT  13.005 1.585 13.125 1.990 ;
        RECT  12.965 1.585 13.005 1.845 ;
        END
        ANTENNAGATEAREA     0.3419 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.605 1.080 17.815 2.315 ;
        RECT  17.295 1.080 17.605 1.290 ;
        RECT  17.355 2.105 17.605 2.315 ;
        RECT  17.295 2.105 17.355 2.585 ;
        RECT  17.035 0.690 17.295 1.290 ;
        RECT  17.035 2.105 17.295 3.045 ;
        END
        ANTENNADIFFAREA     0.8132 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.290 4.265 1.580 ;
        END
        ANTENNAGATEAREA     0.2366 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.290 0.335 2.185 ;
        END
        ANTENNAGATEAREA     0.3783 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 -0.250 17.940 0.250 ;
        RECT  17.545 -0.250 17.805 0.755 ;
        RECT  16.755 -0.250 17.545 0.250 ;
        RECT  16.495 -0.250 16.755 0.405 ;
        RECT  15.195 -0.250 16.495 0.250 ;
        RECT  14.935 -0.250 15.195 0.405 ;
        RECT  12.070 -0.250 14.935 0.250 ;
        RECT  11.810 -0.250 12.070 0.405 ;
        RECT  9.830 -0.250 11.810 0.250 ;
        RECT  9.230 -0.250 9.830 0.405 ;
        RECT  7.615 -0.250 9.230 0.250 ;
        RECT  7.355 -0.250 7.615 0.405 ;
        RECT  6.595 -0.250 7.355 0.250 ;
        RECT  5.995 -0.250 6.595 0.405 ;
        RECT  4.115 -0.250 5.995 0.250 ;
        RECT  3.875 -0.250 4.115 0.405 ;
        RECT  3.515 -0.250 3.875 0.745 ;
        RECT  0.940 -0.250 3.515 0.250 ;
        RECT  0.340 -0.250 0.940 0.405 ;
        RECT  0.000 -0.250 0.340 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 3.440 17.940 3.940 ;
        RECT  17.545 2.615 17.805 3.940 ;
        RECT  16.785 3.440 17.545 3.940 ;
        RECT  16.185 2.955 16.785 3.940 ;
        RECT  14.775 3.440 16.185 3.940 ;
        RECT  14.515 3.285 14.775 3.940 ;
        RECT  12.135 3.440 14.515 3.940 ;
        RECT  11.875 3.285 12.135 3.940 ;
        RECT  10.990 3.440 11.875 3.940 ;
        RECT  10.730 3.285 10.990 3.940 ;
        RECT  9.460 3.440 10.730 3.940 ;
        RECT  9.200 2.660 9.460 3.940 ;
        RECT  6.920 3.440 9.200 3.940 ;
        RECT  6.660 3.285 6.920 3.940 ;
        RECT  1.380 3.440 6.660 3.940 ;
        RECT  0.780 3.285 1.380 3.940 ;
        RECT  0.000 3.440 0.780 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.695 1.495 17.375 1.755 ;
        RECT  16.665 0.695 16.695 1.755 ;
        RECT  16.535 0.695 16.665 2.580 ;
        RECT  15.735 0.695 16.535 0.855 ;
        RECT  16.505 1.495 16.535 2.580 ;
        RECT  16.435 1.495 16.505 1.755 ;
        RECT  15.725 2.420 16.505 2.580 ;
        RECT  16.225 1.035 16.325 1.295 ;
        RECT  16.225 1.955 16.325 2.215 ;
        RECT  16.065 1.035 16.225 2.215 ;
        RECT  15.605 1.725 16.065 1.985 ;
        RECT  15.475 0.695 15.735 1.035 ;
        RECT  15.565 2.420 15.725 2.935 ;
        RECT  13.825 2.775 15.565 2.935 ;
        RECT  13.565 0.840 15.475 1.000 ;
        RECT  15.385 1.215 15.415 1.475 ;
        RECT  15.285 1.215 15.385 2.295 ;
        RECT  15.225 1.215 15.285 2.595 ;
        RECT  15.155 1.215 15.225 1.475 ;
        RECT  15.125 2.035 15.225 2.595 ;
        RECT  14.085 2.435 15.125 2.595 ;
        RECT  14.750 1.180 14.910 2.215 ;
        RECT  13.350 1.180 14.750 1.340 ;
        RECT  14.645 2.055 14.750 2.215 ;
        RECT  13.350 0.470 14.085 0.630 ;
        RECT  13.925 2.005 14.085 2.595 ;
        RECT  13.825 2.005 13.925 2.330 ;
        RECT  12.750 2.170 13.825 2.330 ;
        RECT  13.565 2.775 13.825 3.035 ;
        RECT  13.190 0.470 13.350 1.340 ;
        RECT  12.660 2.515 13.260 2.775 ;
        RECT  12.410 0.470 13.190 0.630 ;
        RECT  12.475 3.060 13.055 3.220 ;
        RECT  12.750 0.810 12.850 1.070 ;
        RECT  12.590 0.810 12.750 2.330 ;
        RECT  10.950 2.605 12.660 2.765 ;
        RECT  11.290 0.925 12.590 1.085 ;
        RECT  12.265 2.065 12.590 2.225 ;
        RECT  12.315 2.945 12.475 3.220 ;
        RECT  12.250 0.470 12.410 0.745 ;
        RECT  10.950 1.265 12.405 1.425 ;
        RECT  10.450 2.945 12.315 3.105 ;
        RECT  12.005 2.015 12.265 2.275 ;
        RECT  11.630 0.585 12.250 0.745 ;
        RECT  11.470 0.470 11.630 0.745 ;
        RECT  10.170 0.470 11.470 0.630 ;
        RECT  11.130 0.810 11.290 1.085 ;
        RECT  10.510 0.810 11.130 0.970 ;
        RECT  10.790 1.150 10.950 2.765 ;
        RECT  10.690 1.150 10.790 1.425 ;
        RECT  10.675 1.870 10.790 2.130 ;
        RECT  10.350 0.810 10.510 1.145 ;
        RECT  10.350 1.385 10.510 1.645 ;
        RECT  10.190 2.945 10.450 3.260 ;
        RECT  7.250 0.985 10.350 1.145 ;
        RECT  10.230 1.485 10.350 1.645 ;
        RECT  10.230 2.605 10.280 2.765 ;
        RECT  10.070 1.485 10.230 2.765 ;
        RECT  9.800 2.945 10.190 3.105 ;
        RECT  10.010 0.470 10.170 0.745 ;
        RECT  9.075 1.485 10.070 1.645 ;
        RECT  10.020 2.605 10.070 2.765 ;
        RECT  9.335 0.585 10.010 0.745 ;
        RECT  9.640 2.210 9.800 3.105 ;
        RECT  8.720 2.210 9.640 2.370 ;
        RECT  9.075 0.585 9.335 0.805 ;
        RECT  4.215 0.585 9.075 0.745 ;
        RECT  8.815 1.325 9.075 1.645 ;
        RECT  8.035 1.485 8.815 1.645 ;
        RECT  8.560 1.925 8.720 3.220 ;
        RECT  8.375 1.925 8.560 2.085 ;
        RECT  7.260 3.060 8.560 3.220 ;
        RECT  7.600 2.720 8.380 2.880 ;
        RECT  8.215 1.825 8.375 2.085 ;
        RECT  8.035 2.350 8.240 2.510 ;
        RECT  7.875 1.485 8.035 2.510 ;
        RECT  7.440 2.605 7.600 2.880 ;
        RECT  6.715 2.605 7.440 2.765 ;
        RECT  7.250 2.265 7.290 2.425 ;
        RECT  7.100 2.945 7.260 3.220 ;
        RECT  7.090 0.935 7.250 2.425 ;
        RECT  6.480 2.945 7.100 3.105 ;
        RECT  6.895 0.935 7.090 1.195 ;
        RECT  7.030 2.265 7.090 2.425 ;
        RECT  6.555 0.925 6.715 2.765 ;
        RECT  5.215 0.925 6.555 1.085 ;
        RECT  5.860 2.395 6.555 2.655 ;
        RECT  6.320 2.945 6.480 3.220 ;
        RECT  1.725 3.060 6.320 3.220 ;
        RECT  5.785 1.865 6.005 2.215 ;
        RECT  5.680 1.275 5.785 2.215 ;
        RECT  5.625 1.275 5.680 2.880 ;
        RECT  4.965 1.275 5.625 1.435 ;
        RECT  5.520 2.055 5.625 2.880 ;
        RECT  2.235 2.720 5.520 2.880 ;
        RECT  4.955 0.925 5.215 1.095 ;
        RECT  4.605 2.040 5.000 2.200 ;
        RECT  4.785 1.275 4.965 1.560 ;
        RECT  4.605 0.925 4.655 1.085 ;
        RECT  4.445 0.925 4.605 2.200 ;
        RECT  4.395 0.925 4.445 1.085 ;
        RECT  4.055 0.585 4.215 1.110 ;
        RECT  3.235 0.950 4.055 1.110 ;
        RECT  3.235 2.040 4.050 2.200 ;
        RECT  3.075 0.930 3.235 2.200 ;
        RECT  2.975 0.930 3.075 1.190 ;
        RECT  2.765 0.470 2.975 0.750 ;
        RECT  2.575 0.930 2.975 1.090 ;
        RECT  1.285 0.470 2.765 0.630 ;
        RECT  2.415 0.810 2.575 1.090 ;
        RECT  1.625 0.810 2.415 0.970 ;
        RECT  2.075 1.150 2.235 2.880 ;
        RECT  1.805 1.150 2.075 1.310 ;
        RECT  1.625 1.575 1.895 1.835 ;
        RECT  1.565 2.120 1.725 3.220 ;
        RECT  1.465 0.810 1.625 1.835 ;
        RECT  1.465 2.120 1.565 2.380 ;
        RECT  1.295 1.575 1.465 1.835 ;
        RECT  1.015 2.120 1.465 2.280 ;
        RECT  1.125 0.470 1.285 0.745 ;
        RECT  1.125 0.970 1.285 1.230 ;
        RECT  0.675 0.585 1.125 0.745 ;
        RECT  1.015 1.070 1.125 1.230 ;
        RECT  0.855 1.070 1.015 2.280 ;
        RECT  0.515 0.585 0.675 2.895 ;
        RECT  0.125 0.835 0.515 1.095 ;
        RECT  0.385 2.735 0.515 2.895 ;
        RECT  0.125 2.735 0.385 2.995 ;
    END
END SDFFSRHQX4

MACRO SDFFSRHQX2
    CLASS CORE ;
    FOREIGN SDFFSRHQX2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.100 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.285 1.580 6.775 1.990 ;
        END
        ANTENNAGATEAREA     0.1911 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.035 1.290 5.395 1.845 ;
        END
        ANTENNAGATEAREA     0.0819 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 1.805 4.515 2.425 ;
        RECT  2.635 2.265 4.355 2.425 ;
        RECT  2.425 2.110 2.635 2.425 ;
        RECT  2.315 2.165 2.425 2.425 ;
        END
        ANTENNAGATEAREA     0.1833 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.755 1.665 12.830 1.925 ;
        RECT  12.570 1.665 12.755 1.990 ;
        RECT  12.545 1.700 12.570 1.990 ;
        RECT  11.955 1.715 12.545 1.875 ;
        RECT  11.795 1.715 11.955 2.055 ;
        RECT  10.795 1.895 11.795 2.055 ;
        END
        ANTENNAGATEAREA     0.2249 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.715 0.695 15.975 1.450 ;
        RECT  15.515 1.290 15.715 1.450 ;
        RECT  15.515 1.925 15.545 2.555 ;
        RECT  15.305 1.290 15.515 2.555 ;
        RECT  15.285 1.955 15.305 2.555 ;
        END
        ANTENNADIFFAREA     0.5668 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.225 1.155 3.635 1.580 ;
        END
        ANTENNAGATEAREA     0.1677 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.290 0.795 1.845 ;
        RECT  0.535 1.585 0.585 1.845 ;
        END
        ANTENNAGATEAREA     0.2314 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.435 -0.250 16.100 0.250 ;
        RECT  15.175 -0.250 15.435 1.090 ;
        RECT  14.835 -0.250 15.175 0.405 ;
        RECT  13.520 -0.250 14.835 0.250 ;
        RECT  13.260 -0.250 13.520 0.405 ;
        RECT  9.065 -0.250 13.260 0.250 ;
        RECT  8.805 -0.250 9.065 0.405 ;
        RECT  5.975 -0.250 8.805 0.250 ;
        RECT  5.715 -0.250 5.975 0.405 ;
        RECT  3.145 -0.250 5.715 0.250 ;
        RECT  2.885 -0.250 3.145 0.405 ;
        RECT  0.935 -0.250 2.885 0.250 ;
        RECT  0.675 -0.250 0.935 0.405 ;
        RECT  0.000 -0.250 0.675 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.945 3.440 16.100 3.940 ;
        RECT  14.885 3.285 15.945 3.940 ;
        RECT  12.935 3.440 14.885 3.940 ;
        RECT  12.675 3.285 12.935 3.940 ;
        RECT  10.515 3.440 12.675 3.940 ;
        RECT  10.255 3.285 10.515 3.940 ;
        RECT  9.565 3.440 10.255 3.940 ;
        RECT  9.305 3.285 9.565 3.940 ;
        RECT  8.315 3.440 9.305 3.940 ;
        RECT  8.055 3.285 8.315 3.940 ;
        RECT  6.005 3.440 8.055 3.940 ;
        RECT  5.745 3.285 6.005 3.940 ;
        RECT  3.775 3.440 5.745 3.940 ;
        RECT  3.515 3.285 3.775 3.940 ;
        RECT  1.405 3.440 3.515 3.940 ;
        RECT  0.725 3.285 1.405 3.940 ;
        RECT  0.465 2.890 0.725 3.940 ;
        RECT  0.000 3.440 0.465 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.975 1.580 15.105 1.840 ;
        RECT  14.815 0.675 14.975 3.085 ;
        RECT  14.095 0.675 14.815 0.835 ;
        RECT  12.200 2.925 14.815 3.085 ;
        RECT  14.425 2.465 14.635 2.725 ;
        RECT  14.425 1.035 14.525 1.295 ;
        RECT  14.265 1.035 14.425 2.725 ;
        RECT  14.005 1.495 14.265 1.755 ;
        RECT  13.835 0.525 14.095 0.835 ;
        RECT  13.785 1.015 14.005 1.275 ;
        RECT  12.320 0.675 13.835 0.835 ;
        RECT  13.685 1.015 13.785 2.450 ;
        RECT  13.625 1.015 13.685 2.745 ;
        RECT  13.525 2.190 13.625 2.745 ;
        RECT  12.540 2.585 13.525 2.745 ;
        RECT  13.255 2.145 13.305 2.405 ;
        RECT  13.095 1.235 13.255 2.405 ;
        RECT  11.880 1.235 13.095 1.395 ;
        RECT  13.045 2.145 13.095 2.405 ;
        RECT  12.395 2.265 12.540 2.745 ;
        RECT  12.380 2.165 12.395 2.745 ;
        RECT  12.135 2.165 12.380 2.425 ;
        RECT  12.060 0.675 12.320 1.055 ;
        RECT  12.040 2.655 12.200 3.085 ;
        RECT  10.610 2.265 12.135 2.425 ;
        RECT  11.940 2.655 12.040 2.915 ;
        RECT  11.720 0.470 11.880 1.395 ;
        RECT  9.405 0.470 11.720 0.630 ;
        RECT  11.205 2.605 11.465 2.885 ;
        RECT  11.255 0.810 11.415 1.715 ;
        RECT  11.025 3.065 11.365 3.225 ;
        RECT  9.745 0.810 11.255 0.970 ;
        RECT  10.610 1.555 11.255 1.715 ;
        RECT  10.115 2.605 11.205 2.765 ;
        RECT  10.130 1.205 11.075 1.365 ;
        RECT  10.865 2.945 11.025 3.225 ;
        RECT  9.025 2.945 10.865 3.105 ;
        RECT  10.450 1.555 10.610 2.425 ;
        RECT  10.315 2.265 10.450 2.425 ;
        RECT  9.970 1.205 10.130 1.425 ;
        RECT  9.955 2.185 10.115 2.765 ;
        RECT  9.470 1.265 9.970 1.425 ;
        RECT  9.470 2.185 9.955 2.345 ;
        RECT  9.585 0.810 9.745 1.085 ;
        RECT  8.285 0.925 9.585 1.085 ;
        RECT  9.310 1.265 9.470 2.345 ;
        RECT  9.245 0.470 9.405 0.745 ;
        RECT  9.075 1.935 9.310 2.195 ;
        RECT  8.625 0.585 9.245 0.745 ;
        RECT  8.895 1.455 9.130 1.715 ;
        RECT  8.765 2.945 9.025 3.205 ;
        RECT  8.735 1.455 8.895 2.760 ;
        RECT  7.235 2.945 8.765 3.105 ;
        RECT  8.565 2.500 8.735 2.760 ;
        RECT  8.465 0.470 8.625 0.745 ;
        RECT  7.555 2.600 8.565 2.760 ;
        RECT  6.315 0.470 8.465 0.630 ;
        RECT  8.125 0.810 8.285 1.085 ;
        RECT  6.655 0.810 8.125 0.970 ;
        RECT  7.765 1.150 7.945 1.310 ;
        RECT  7.605 1.150 7.765 2.270 ;
        RECT  7.555 2.110 7.605 2.270 ;
        RECT  7.395 2.110 7.555 2.760 ;
        RECT  7.215 1.445 7.265 1.705 ;
        RECT  7.215 2.945 7.235 3.210 ;
        RECT  7.055 1.445 7.215 3.210 ;
        RECT  7.005 1.445 7.055 1.705 ;
        RECT  6.345 3.050 7.055 3.210 ;
        RECT  6.715 2.555 6.875 2.870 ;
        RECT  5.735 2.555 6.715 2.715 ;
        RECT  6.495 0.810 6.655 1.110 ;
        RECT  6.075 0.950 6.495 1.110 ;
        RECT  6.185 2.945 6.345 3.210 ;
        RECT  6.155 0.470 6.315 0.745 ;
        RECT  3.045 2.945 6.185 3.105 ;
        RECT  5.535 0.585 6.155 0.745 ;
        RECT  5.915 0.950 6.075 2.255 ;
        RECT  5.575 0.925 5.735 2.715 ;
        RECT  5.195 0.925 5.575 1.085 ;
        RECT  5.195 2.505 5.575 2.715 ;
        RECT  5.375 0.475 5.535 0.745 ;
        RECT  4.855 2.115 5.390 2.275 ;
        RECT  3.485 0.475 5.375 0.635 ;
        RECT  5.035 0.815 5.195 1.085 ;
        RECT  5.035 2.505 5.195 2.765 ;
        RECT  4.225 0.815 5.035 0.975 ;
        RECT  4.695 1.335 4.855 2.765 ;
        RECT  4.315 1.335 4.695 1.495 ;
        RECT  2.705 2.605 4.695 2.765 ;
        RECT  4.155 1.155 4.315 1.495 ;
        RECT  3.975 1.925 4.175 2.085 ;
        RECT  3.815 0.815 3.975 2.085 ;
        RECT  3.715 0.815 3.815 0.975 ;
        RECT  3.325 0.475 3.485 0.970 ;
        RECT  2.975 0.810 3.325 0.970 ;
        RECT  2.975 1.925 3.225 2.085 ;
        RECT  2.885 2.945 3.045 3.220 ;
        RECT  2.815 0.810 2.975 2.085 ;
        RECT  1.765 3.060 2.885 3.220 ;
        RECT  2.555 0.810 2.815 1.075 ;
        RECT  2.445 2.605 2.705 2.880 ;
        RECT  1.705 0.810 2.555 0.970 ;
        RECT  2.135 2.605 2.445 2.765 ;
        RECT  2.135 1.150 2.305 1.310 ;
        RECT  1.310 0.460 2.145 0.620 ;
        RECT  1.975 1.150 2.135 2.765 ;
        RECT  1.605 2.070 1.765 3.220 ;
        RECT  1.545 0.810 1.705 1.845 ;
        RECT  1.505 2.070 1.605 2.670 ;
        RECT  1.335 1.585 1.545 1.845 ;
        RECT  1.135 2.070 1.505 2.230 ;
        RECT  1.135 1.035 1.365 1.295 ;
        RECT  1.150 0.460 1.310 0.750 ;
        RECT  0.385 0.590 1.150 0.750 ;
        RECT  0.975 1.035 1.135 2.230 ;
        RECT  0.285 0.590 0.385 1.290 ;
        RECT  0.285 2.025 0.385 2.285 ;
        RECT  0.225 0.590 0.285 2.285 ;
        RECT  0.125 1.030 0.225 2.285 ;
    END
END SDFFSRHQX2

MACRO SDFFSRHQX1
    CLASS CORE ;
    FOREIGN SDFFSRHQX1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.180 BY 3.690 ;
    SYMMETRY X Y ;
    SITE TSM13SITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.975 1.330 6.315 2.150 ;
        END
        ANTENNAGATEAREA     0.1365 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.290 5.040 1.845 ;
        RECT  4.725 1.290 4.820 1.580 ;
        END
        ANTENNAGATEAREA     0.0494 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 2.100 4.235 2.540 ;
        RECT  3.135 2.380 4.075 2.540 ;
        RECT  2.975 1.290 3.135 2.540 ;
        RECT  2.885 1.290 2.975 1.580 ;
        RECT  2.355 2.380 2.975 2.540 ;
        RECT  2.195 2.165 2.355 2.540 ;
        END
        ANTENNAGATEAREA     0.1261 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.880 1.635 12.140 1.895 ;
        RECT  11.810 1.685 11.880 1.895 ;
        RECT  10.475 1.685 11.810 1.845 ;
        RECT  10.245 1.300 10.475 1.990 ;
        END
        ANTENNAGATEAREA     0.1404 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.975 1.290 15.055 2.175 ;
        RECT  14.715 1.035 14.975 2.555 ;
        END
        ANTENNADIFFAREA     0.3944 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.315 1.290 3.555 1.860 ;
        END
        ANTENNAGATEAREA     0.0962 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.125 1.180 0.435 1.845 ;
        END
        ANTENNAGATEAREA     0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.425 -0.250 15.180 0.250 ;
        RECT  14.165 -0.250 14.425 0.405 ;
        RECT  12.825 -0.250 14.165 0.250 ;
        RECT  12.565 -0.250 12.825 0.405 ;
        RECT  10.305 -0.250 12.565 0.250 ;
        RECT  10.045 -0.250 10.305 0.405 ;
        RECT  8.700 -0.250 10.045 0.250 ;
        RECT  8.440 -0.250 8.700 0.405 ;
        RECT  5.045 -0.250 8.440 0.250 ;
        RECT  4.785 -0.250 5.045 0.405 ;
        RECT  3.205 -0.250 4.785 0.250 ;
        RECT  2.945 -0.250 3.205 0.405 ;
        RECT  0.895 -0.250 2.945 0.250 ;
        RECT  0.635 -0.250 0.895 0.405 ;
        RECT  0.000 -0.250 0.635 0.250 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.425 3.440 15.180 3.940 ;
        RECT  13.825 2.880 14.425 3.940 ;
        RECT  12.435 3.440 13.825 3.940 ;
        RECT  12.175 3.285 12.435 3.940 ;
        RECT  9.155 3.440 12.175 3.940 ;
        RECT  8.895 3.285 9.155 3.940 ;
        RECT  7.755 3.440 8.895 3.940 ;
        RECT  7.495 3.285 7.755 3.940 ;
        RECT  5.635 3.440 7.495 3.940 ;
        RECT  5.375 3.285 5.635 3.940 ;
        RECT  1.235 3.440 5.375 3.940 ;
        RECT  0.635 3.285 1.235 3.940 ;
        RECT  0.000 3.440 0.635 3.940 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.205 0.625 14.365 2.695 ;
        RECT  13.515 0.625 14.205 0.785 ;
        RECT  14.105 1.515 14.205 1.775 ;
        RECT  12.945 2.535 14.205 2.695 ;
        RECT  13.895 1.035 13.995 1.295 ;
        RECT  13.895 1.955 13.995 2.215 ;
        RECT  13.735 1.035 13.895 2.215 ;
        RECT  13.535 1.445 13.735 1.705 ;
        RECT  13.255 0.525 13.515 0.785 ;
        RECT  13.215 0.965 13.315 1.225 ;
        RECT  13.215 1.755 13.315 2.015 ;
        RECT  11.630 0.625 13.255 0.785 ;
        RECT  13.055 0.965 13.215 2.355 ;
        RECT  11.305 2.195 13.055 2.355 ;
        RECT  12.685 2.535 12.945 3.155 ;
        RECT  12.735 1.755 12.835 2.015 ;
        RECT  12.575 1.295 12.735 2.015 ;
        RECT  11.645 2.535 12.685 2.695 ;
        RECT  11.190 1.295 12.575 1.455 ;
        RECT  11.485 2.535 11.645 2.810 ;
        RECT  11.470 0.625 11.630 1.065 ;
        RECT  11.370 0.805 11.470 1.065 ;
        RECT  11.145 2.195 11.305 2.760 ;
        RECT  11.030 0.455 11.190 1.455 ;
        RECT  8.555 2.600 11.1